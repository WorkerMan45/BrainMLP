// hps.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module hps (
		output wire [15:0] address_external_connection_export,         //       address_external_connection.export
		input  wire        clk_clk,                                    //                               clk.clk
		output wire        clock_in_external_connection_export,        //      clock_in_external_connection.export
		output wire [31:0] din_external_connection_export,             //           din_external_connection.export
		input  wire [31:0] dout_external_connection_export,            //          dout_external_connection.export
		input  wire [7:0]  enableregions_external_connection_in_port,  // enableregions_external_connection.in_port
		output wire [7:0]  enableregions_external_connection_out_port, //                                  .out_port
		output wire        hps_io_hps_io_emac1_inst_TX_CLK,            //                            hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,              //                                  .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,              //                                  .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,              //                                  .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,              //                                  .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,              //                                  .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,              //                                  .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,               //                                  .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL,            //                                  .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL,            //                                  .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK,            //                                  .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,              //                                  .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,              //                                  .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,              //                                  .hps_io_emac1_inst_RXD3
		inout  wire        hps_io_hps_io_sdio_inst_CMD,                //                                  .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,                 //                                  .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,                 //                                  .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,                //                                  .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,                 //                                  .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,                 //                                  .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,                 //                                  .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,                 //                                  .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,                 //                                  .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,                 //                                  .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,                 //                                  .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,                 //                                  .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,                 //                                  .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,                 //                                  .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,                //                                  .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,                //                                  .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,                //                                  .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,                //                                  .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,                //                                  .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,                //                                  .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_gpio_inst_GPIO35,             //                                  .hps_io_gpio_inst_GPIO35
		input  wire [31:0] layer1_external_connection_in_port,         //        layer1_external_connection.in_port
		output wire [31:0] layer1_external_connection_out_port,        //                                  .out_port
		input  wire [31:0] layer2_external_connection_in_port,         //        layer2_external_connection.in_port
		output wire [31:0] layer2_external_connection_out_port,        //                                  .out_port
		input  wire [31:0] layer3_external_connection_in_port,         //        layer3_external_connection.in_port
		output wire [31:0] layer3_external_connection_out_port,        //                                  .out_port
		output wire [14:0] memory_mem_a,                               //                            memory.mem_a
		output wire [2:0]  memory_mem_ba,                              //                                  .mem_ba
		output wire        memory_mem_ck,                              //                                  .mem_ck
		output wire        memory_mem_ck_n,                            //                                  .mem_ck_n
		output wire        memory_mem_cke,                             //                                  .mem_cke
		output wire        memory_mem_cs_n,                            //                                  .mem_cs_n
		output wire        memory_mem_ras_n,                           //                                  .mem_ras_n
		output wire        memory_mem_cas_n,                           //                                  .mem_cas_n
		output wire        memory_mem_we_n,                            //                                  .mem_we_n
		output wire        memory_mem_reset_n,                         //                                  .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                              //                                  .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                             //                                  .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                           //                                  .mem_dqs_n
		output wire        memory_mem_odt,                             //                                  .mem_odt
		output wire [3:0]  memory_mem_dm,                              //                                  .mem_dm
		input  wire        memory_oct_rzqin,                           //                                  .oct_rzqin
		output wire        read_external_connection_export,            //          read_external_connection.export
		output wire        reset_in_external_connection_export,        //      reset_in_external_connection.export
		output wire        write_external_connection_export            //         write_external_connection.export
	);

	wire         hps_0_h2f_reset_reset;                         // hps_0:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;               // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                 // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                 // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                 // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                   // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;               // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                 // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;               // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;               // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                  // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;               // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;               // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;               // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                 // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                 // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                  // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;               // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_write_s1_chipselect;         // mm_interconnect_0:Write_s1_chipselect -> Write:chipselect
	wire  [31:0] mm_interconnect_0_write_s1_readdata;           // Write:readdata -> mm_interconnect_0:Write_s1_readdata
	wire   [1:0] mm_interconnect_0_write_s1_address;            // mm_interconnect_0:Write_s1_address -> Write:address
	wire         mm_interconnect_0_write_s1_write;              // mm_interconnect_0:Write_s1_write -> Write:write_n
	wire  [31:0] mm_interconnect_0_write_s1_writedata;          // mm_interconnect_0:Write_s1_writedata -> Write:writedata
	wire         mm_interconnect_0_address_s1_chipselect;       // mm_interconnect_0:Address_s1_chipselect -> Address:chipselect
	wire  [31:0] mm_interconnect_0_address_s1_readdata;         // Address:readdata -> mm_interconnect_0:Address_s1_readdata
	wire   [1:0] mm_interconnect_0_address_s1_address;          // mm_interconnect_0:Address_s1_address -> Address:address
	wire         mm_interconnect_0_address_s1_write;            // mm_interconnect_0:Address_s1_write -> Address:write_n
	wire  [31:0] mm_interconnect_0_address_s1_writedata;        // mm_interconnect_0:Address_s1_writedata -> Address:writedata
	wire         mm_interconnect_0_din_s1_chipselect;           // mm_interconnect_0:Din_s1_chipselect -> Din:chipselect
	wire  [31:0] mm_interconnect_0_din_s1_readdata;             // Din:readdata -> mm_interconnect_0:Din_s1_readdata
	wire   [1:0] mm_interconnect_0_din_s1_address;              // mm_interconnect_0:Din_s1_address -> Din:address
	wire         mm_interconnect_0_din_s1_write;                // mm_interconnect_0:Din_s1_write -> Din:write_n
	wire  [31:0] mm_interconnect_0_din_s1_writedata;            // mm_interconnect_0:Din_s1_writedata -> Din:writedata
	wire  [31:0] mm_interconnect_0_dout_s1_readdata;            // Dout:readdata -> mm_interconnect_0:Dout_s1_readdata
	wire   [1:0] mm_interconnect_0_dout_s1_address;             // mm_interconnect_0:Dout_s1_address -> Dout:address
	wire         mm_interconnect_0_reset_in_s1_chipselect;      // mm_interconnect_0:Reset_In_s1_chipselect -> Reset_In:chipselect
	wire  [31:0] mm_interconnect_0_reset_in_s1_readdata;        // Reset_In:readdata -> mm_interconnect_0:Reset_In_s1_readdata
	wire   [1:0] mm_interconnect_0_reset_in_s1_address;         // mm_interconnect_0:Reset_In_s1_address -> Reset_In:address
	wire         mm_interconnect_0_reset_in_s1_write;           // mm_interconnect_0:Reset_In_s1_write -> Reset_In:write_n
	wire  [31:0] mm_interconnect_0_reset_in_s1_writedata;       // mm_interconnect_0:Reset_In_s1_writedata -> Reset_In:writedata
	wire         mm_interconnect_0_enableregions_s1_chipselect; // mm_interconnect_0:EnableRegions_s1_chipselect -> EnableRegions:chipselect
	wire  [31:0] mm_interconnect_0_enableregions_s1_readdata;   // EnableRegions:readdata -> mm_interconnect_0:EnableRegions_s1_readdata
	wire   [1:0] mm_interconnect_0_enableregions_s1_address;    // mm_interconnect_0:EnableRegions_s1_address -> EnableRegions:address
	wire         mm_interconnect_0_enableregions_s1_write;      // mm_interconnect_0:EnableRegions_s1_write -> EnableRegions:write_n
	wire  [31:0] mm_interconnect_0_enableregions_s1_writedata;  // mm_interconnect_0:EnableRegions_s1_writedata -> EnableRegions:writedata
	wire         mm_interconnect_0_layer1_s1_chipselect;        // mm_interconnect_0:Layer1_s1_chipselect -> Layer1:chipselect
	wire  [31:0] mm_interconnect_0_layer1_s1_readdata;          // Layer1:readdata -> mm_interconnect_0:Layer1_s1_readdata
	wire   [1:0] mm_interconnect_0_layer1_s1_address;           // mm_interconnect_0:Layer1_s1_address -> Layer1:address
	wire         mm_interconnect_0_layer1_s1_write;             // mm_interconnect_0:Layer1_s1_write -> Layer1:write_n
	wire  [31:0] mm_interconnect_0_layer1_s1_writedata;         // mm_interconnect_0:Layer1_s1_writedata -> Layer1:writedata
	wire         mm_interconnect_0_layer2_s1_chipselect;        // mm_interconnect_0:Layer2_s1_chipselect -> Layer2:chipselect
	wire  [31:0] mm_interconnect_0_layer2_s1_readdata;          // Layer2:readdata -> mm_interconnect_0:Layer2_s1_readdata
	wire   [1:0] mm_interconnect_0_layer2_s1_address;           // mm_interconnect_0:Layer2_s1_address -> Layer2:address
	wire         mm_interconnect_0_layer2_s1_write;             // mm_interconnect_0:Layer2_s1_write -> Layer2:write_n
	wire  [31:0] mm_interconnect_0_layer2_s1_writedata;         // mm_interconnect_0:Layer2_s1_writedata -> Layer2:writedata
	wire         mm_interconnect_0_layer3_s1_chipselect;        // mm_interconnect_0:Layer3_s1_chipselect -> Layer3:chipselect
	wire  [31:0] mm_interconnect_0_layer3_s1_readdata;          // Layer3:readdata -> mm_interconnect_0:Layer3_s1_readdata
	wire   [1:0] mm_interconnect_0_layer3_s1_address;           // mm_interconnect_0:Layer3_s1_address -> Layer3:address
	wire         mm_interconnect_0_layer3_s1_write;             // mm_interconnect_0:Layer3_s1_write -> Layer3:write_n
	wire  [31:0] mm_interconnect_0_layer3_s1_writedata;         // mm_interconnect_0:Layer3_s1_writedata -> Layer3:writedata
	wire         mm_interconnect_0_clock_in_s1_chipselect;      // mm_interconnect_0:Clock_In_s1_chipselect -> Clock_In:chipselect
	wire  [31:0] mm_interconnect_0_clock_in_s1_readdata;        // Clock_In:readdata -> mm_interconnect_0:Clock_In_s1_readdata
	wire   [1:0] mm_interconnect_0_clock_in_s1_address;         // mm_interconnect_0:Clock_In_s1_address -> Clock_In:address
	wire         mm_interconnect_0_clock_in_s1_write;           // mm_interconnect_0:Clock_In_s1_write -> Clock_In:write_n
	wire  [31:0] mm_interconnect_0_clock_in_s1_writedata;       // mm_interconnect_0:Clock_In_s1_writedata -> Clock_In:writedata
	wire         mm_interconnect_0_read_s1_chipselect;          // mm_interconnect_0:Read_s1_chipselect -> Read:chipselect
	wire  [31:0] mm_interconnect_0_read_s1_readdata;            // Read:readdata -> mm_interconnect_0:Read_s1_readdata
	wire   [1:0] mm_interconnect_0_read_s1_address;             // mm_interconnect_0:Read_s1_address -> Read:address
	wire         mm_interconnect_0_read_s1_write;               // mm_interconnect_0:Read_s1_write -> Read:write_n
	wire  [31:0] mm_interconnect_0_read_s1_writedata;           // mm_interconnect_0:Read_s1_writedata -> Read:writedata
	wire         rst_controller_reset_out_reset;                // rst_controller:reset_out -> [Address:reset_n, Clock_In:reset_n, Din:reset_n, Dout:reset_n, EnableRegions:reset_n, Layer1:reset_n, Layer2:reset_n, Layer3:reset_n, Read:reset_n, Reset_In:reset_n, Write:reset_n, mm_interconnect_0:Write_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;            // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	hps_Address address (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_address_s1_readdata),   //                    .readdata
		.out_port   (address_external_connection_export)       // external_connection.export
	);

	hps_Clock_In clock_in (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_clock_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_clock_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_clock_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_clock_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_clock_in_s1_readdata),   //                    .readdata
		.out_port   (clock_in_external_connection_export)       // external_connection.export
	);

	hps_Din din (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_din_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_din_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_din_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_din_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_din_s1_readdata),   //                    .readdata
		.out_port   (din_external_connection_export)       // external_connection.export
	);

	hps_Dout dout (
		.clk      (clk_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address  (mm_interconnect_0_dout_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_dout_s1_readdata), //                    .readdata
		.in_port  (dout_external_connection_export)     // external_connection.export
	);

	hps_EnableRegions enableregions (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_enableregions_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_enableregions_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_enableregions_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_enableregions_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_enableregions_s1_readdata),   //                    .readdata
		.in_port    (enableregions_external_connection_in_port),     // external_connection.export
		.out_port   (enableregions_external_connection_out_port)     //                    .export
	);

	hps_Layer1 layer1 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_layer1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_layer1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_layer1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_layer1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_layer1_s1_readdata),   //                    .readdata
		.in_port    (layer1_external_connection_in_port),     // external_connection.export
		.out_port   (layer1_external_connection_out_port)     //                    .export
	);

	hps_Layer1 layer2 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_layer2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_layer2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_layer2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_layer2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_layer2_s1_readdata),   //                    .readdata
		.in_port    (layer2_external_connection_in_port),     // external_connection.export
		.out_port   (layer2_external_connection_out_port)     //                    .export
	);

	hps_Layer1 layer3 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_layer3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_layer3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_layer3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_layer3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_layer3_s1_readdata),   //                    .readdata
		.in_port    (layer3_external_connection_in_port),     // external_connection.export
		.out_port   (layer3_external_connection_out_port)     //                    .export
	);

	hps_Clock_In read (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_read_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_read_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_read_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_read_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_read_s1_readdata),   //                    .readdata
		.out_port   (read_external_connection_export)       // external_connection.export
	);

	hps_Clock_In reset_in (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_reset_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_in_s1_readdata),   //                    .readdata
		.out_port   (reset_in_external_connection_export)       // external_connection.export
	);

	hps_Clock_In write (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_write_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_write_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_write_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_write_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_write_s1_readdata),   //                    .readdata
		.out_port   (write_external_connection_export)       // external_connection.export
	);

	hps_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                    //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                   //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                   //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                 //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                  //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                 //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                 //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),              //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                   //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                  //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                  //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                   //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready)   //                  .rready
	);

	hps_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                  //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                 //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),               //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),               //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),               //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),               //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                   //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                 //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                 //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                 //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                   //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                 //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                  //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                 //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),               //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),               //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),               //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),               //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                   //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                 //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                 //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                 //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                       //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),            // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.Write_reset_reset_bridge_in_reset_reset                             (rst_controller_reset_out_reset),                //                             Write_reset_reset_bridge_in_reset.reset
		.Address_s1_address                                                  (mm_interconnect_0_address_s1_address),          //                                                    Address_s1.address
		.Address_s1_write                                                    (mm_interconnect_0_address_s1_write),            //                                                              .write
		.Address_s1_readdata                                                 (mm_interconnect_0_address_s1_readdata),         //                                                              .readdata
		.Address_s1_writedata                                                (mm_interconnect_0_address_s1_writedata),        //                                                              .writedata
		.Address_s1_chipselect                                               (mm_interconnect_0_address_s1_chipselect),       //                                                              .chipselect
		.Clock_In_s1_address                                                 (mm_interconnect_0_clock_in_s1_address),         //                                                   Clock_In_s1.address
		.Clock_In_s1_write                                                   (mm_interconnect_0_clock_in_s1_write),           //                                                              .write
		.Clock_In_s1_readdata                                                (mm_interconnect_0_clock_in_s1_readdata),        //                                                              .readdata
		.Clock_In_s1_writedata                                               (mm_interconnect_0_clock_in_s1_writedata),       //                                                              .writedata
		.Clock_In_s1_chipselect                                              (mm_interconnect_0_clock_in_s1_chipselect),      //                                                              .chipselect
		.Din_s1_address                                                      (mm_interconnect_0_din_s1_address),              //                                                        Din_s1.address
		.Din_s1_write                                                        (mm_interconnect_0_din_s1_write),                //                                                              .write
		.Din_s1_readdata                                                     (mm_interconnect_0_din_s1_readdata),             //                                                              .readdata
		.Din_s1_writedata                                                    (mm_interconnect_0_din_s1_writedata),            //                                                              .writedata
		.Din_s1_chipselect                                                   (mm_interconnect_0_din_s1_chipselect),           //                                                              .chipselect
		.Dout_s1_address                                                     (mm_interconnect_0_dout_s1_address),             //                                                       Dout_s1.address
		.Dout_s1_readdata                                                    (mm_interconnect_0_dout_s1_readdata),            //                                                              .readdata
		.EnableRegions_s1_address                                            (mm_interconnect_0_enableregions_s1_address),    //                                              EnableRegions_s1.address
		.EnableRegions_s1_write                                              (mm_interconnect_0_enableregions_s1_write),      //                                                              .write
		.EnableRegions_s1_readdata                                           (mm_interconnect_0_enableregions_s1_readdata),   //                                                              .readdata
		.EnableRegions_s1_writedata                                          (mm_interconnect_0_enableregions_s1_writedata),  //                                                              .writedata
		.EnableRegions_s1_chipselect                                         (mm_interconnect_0_enableregions_s1_chipselect), //                                                              .chipselect
		.Layer1_s1_address                                                   (mm_interconnect_0_layer1_s1_address),           //                                                     Layer1_s1.address
		.Layer1_s1_write                                                     (mm_interconnect_0_layer1_s1_write),             //                                                              .write
		.Layer1_s1_readdata                                                  (mm_interconnect_0_layer1_s1_readdata),          //                                                              .readdata
		.Layer1_s1_writedata                                                 (mm_interconnect_0_layer1_s1_writedata),         //                                                              .writedata
		.Layer1_s1_chipselect                                                (mm_interconnect_0_layer1_s1_chipselect),        //                                                              .chipselect
		.Layer2_s1_address                                                   (mm_interconnect_0_layer2_s1_address),           //                                                     Layer2_s1.address
		.Layer2_s1_write                                                     (mm_interconnect_0_layer2_s1_write),             //                                                              .write
		.Layer2_s1_readdata                                                  (mm_interconnect_0_layer2_s1_readdata),          //                                                              .readdata
		.Layer2_s1_writedata                                                 (mm_interconnect_0_layer2_s1_writedata),         //                                                              .writedata
		.Layer2_s1_chipselect                                                (mm_interconnect_0_layer2_s1_chipselect),        //                                                              .chipselect
		.Layer3_s1_address                                                   (mm_interconnect_0_layer3_s1_address),           //                                                     Layer3_s1.address
		.Layer3_s1_write                                                     (mm_interconnect_0_layer3_s1_write),             //                                                              .write
		.Layer3_s1_readdata                                                  (mm_interconnect_0_layer3_s1_readdata),          //                                                              .readdata
		.Layer3_s1_writedata                                                 (mm_interconnect_0_layer3_s1_writedata),         //                                                              .writedata
		.Layer3_s1_chipselect                                                (mm_interconnect_0_layer3_s1_chipselect),        //                                                              .chipselect
		.Read_s1_address                                                     (mm_interconnect_0_read_s1_address),             //                                                       Read_s1.address
		.Read_s1_write                                                       (mm_interconnect_0_read_s1_write),               //                                                              .write
		.Read_s1_readdata                                                    (mm_interconnect_0_read_s1_readdata),            //                                                              .readdata
		.Read_s1_writedata                                                   (mm_interconnect_0_read_s1_writedata),           //                                                              .writedata
		.Read_s1_chipselect                                                  (mm_interconnect_0_read_s1_chipselect),          //                                                              .chipselect
		.Reset_In_s1_address                                                 (mm_interconnect_0_reset_in_s1_address),         //                                                   Reset_In_s1.address
		.Reset_In_s1_write                                                   (mm_interconnect_0_reset_in_s1_write),           //                                                              .write
		.Reset_In_s1_readdata                                                (mm_interconnect_0_reset_in_s1_readdata),        //                                                              .readdata
		.Reset_In_s1_writedata                                               (mm_interconnect_0_reset_in_s1_writedata),       //                                                              .writedata
		.Reset_In_s1_chipselect                                              (mm_interconnect_0_reset_in_s1_chipselect),      //                                                              .chipselect
		.Write_s1_address                                                    (mm_interconnect_0_write_s1_address),            //                                                      Write_s1.address
		.Write_s1_write                                                      (mm_interconnect_0_write_s1_write),              //                                                              .write
		.Write_s1_readdata                                                   (mm_interconnect_0_write_s1_readdata),           //                                                              .readdata
		.Write_s1_writedata                                                  (mm_interconnect_0_write_s1_writedata),          //                                                              .writedata
		.Write_s1_chipselect                                                 (mm_interconnect_0_write_s1_chipselect)          //                                                              .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
