library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity grebal_vga8_20x20 is
port (
	clk, en : in std_logic;
	addr : in unsigned(15 downto 0);
	data : out unsigned(27 downto 0));
end grebal_vga8_20x20;

architecture imp of grebal_vga8_20x20 is
	type rom_type is array (0 to 50297) of unsigned(27 downto 0); -- unused[3]; is_background[1]; R[8]; G[8]; B[8]
	constant ROM : rom_type :=
	(
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110011111100111111001","0000111110001111100011111000","0000111110001111100011111000","0000111111101111111011111110","0000111101011111010111110101","0000111011111110111111101111","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100111111001111110011","0000111111111111111111111111","0000111100001111000011110000","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000110010011100100111001001","0000101001011010010110100101","0000011101100111011001110110","0000001101100011011000110110","0000000111000001110000011100","0001000000000000000000000000","0001000000000000000000000000","0000000111100001111000011110","0000011010100110101001101010","0000101011001010110010101100","0000111100011111000111110001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110011111100111111001","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111100001111000011110000","0000111100011111000111110001","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000101110011011100110111001","0000101100001011000010110000","0000100101111001011110010111","0000100110001001100010011000","0000100100101001001010010010","0000101011101010111010101110","0000101111001011110010111100","0000110011111100111111001111","0000111011001110110011101100","0000111100011111000111110001","0000111110001111100011111000","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101011111010111110101","0000111111101111111011111110","0000111101111111011111110111","0000111101011111010111110101","0000111111011111110111111101","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111100101111001011110010","0000111100101111001011110010","0000111110011111100111111001","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111101011111010111110101","0000111110011111100111111001","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111010101110101011101010","0000110011011100110111001101","0000100110011001100110011001","0000010011000100110001001100","0000000010100000101000001010","0000001000110010001100100011","0000100001111000011110000111","0000100001011000010110000101","0000100100101001001010010010","0000101001001010010010100100","0000110010111100101111001011","0000110101011101010111010101","0000100110001001100010011000","0000011010000110100001101000","0000001010010010100100101001","0000100100111001001110010011","0000111000011110000111100001","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111100001111000011110000","0000111111101111111011111110","0000111101011111010111110101","0000111111011111110111111101","0000101110011011100110111001","0000011000110110001101100011","0001000000000000000000000000","0000000110010001100100011001","0000001101100011011000110110","0000001100010011000100110001","0000001001000010010000100100","0000000100000001000000010000","0000001000100010001000100010","0000000011010000110100001101","0001000000000000000000000000","0001000000000000000000000000","0000000111010001110100011101","0000010001100100011001000110","0000100011111000111110001111","0000101111001011110010111100","0000110011111100111111001111","0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111100101111001011110010","0000111100001111000011110000","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111111101111111011111110","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000110111101101111011011110","0000101001101010011010100110","0000001101100011011000110110","0000001000010010000100100001","0000001101100011011000110110","0000010001000100010001000100","0000010000010100000101000001","0000011001000110010001100100","0000100110101001101010011010","0000100101001001010010010100","0000101001111010011110100111","0000101101001011010010110100","0000100000001000000010000000","0000101000101010001010100010","0000110011111100111111001111","0000110101011101010111010101","0000101100111011001110110011","0000010011100100111001001110","0000001111110011111100111111","0000110101001101010011010100","0000111101001111010011110100","0000111111111111111111111111","0000111100011111000111110001","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111101101111011011110110","0000110101101101011011010110","0000010101000101010001010100","0001000000000000000000000000","0000001000110010001100100011","0000100000001000000010000000","0000101100111011001110110011","0000101100101011001010110010","0000101011001010110010101100","0000101101101011011010110110","0000100110011001100110011001","0000100010101000101010001010","0000011101110111011101110111","0000100000001000000010000000","0000100011001000110010001100","0000011011000110110001101100","0000011101010111010101110101","0000011011110110111101101111","0000010000000100000001000000","0000001011000010110000101100","0000010001000100010001000100","0000011000110110001101100011","0000100111101001111010011110","0000110011101100111011001110","0000110001111100011111000111","0000110000001100000011000000","0000111010001110100011101000","0000111011011110110111101101","0000111000101110001011100010","0000111111111111111111111111","0000111101101111011011110110","0000111101001111010011110100","0000111111011111110111111101","0000111100101111001011110010","0000111111011111110111111101","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111011011110110111101101","0000111101001111010011110100","0000111110011111100111111001","0000111101111111011111110111","0000111100101111001011110010","0000111101001111010011110100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101011111010111110101","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101111111011111110111","0000111110001111100011111000","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000110011111100111111001111","0000011110000111100001111000","0000001010010010100100101001","0000001100100011001000110010","0000011111100111111001111110","0000100100111001001110010011","0000010101110101011101010111","0000011111100111111001111110","0000011100010111000101110001","0000011101000111010001110100","0000011101010111010101110101","0000100100001001000010010000","0000100010001000100010001000","0000110100111101001111010011","0000110000001100000011000000","0000110001111100011111000111","0000101010101010101010101010","0000101010101010101010101010","0000101000011010000110100001","0000100000111000001110000011","0000010111100101111001011110","0001000000000000000000000000","0000110101111101011111010111","0000111111111111111111111111","0000111111001111110011111100","0000111100111111001111110011","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000101010111010101110101011","0001000000000000000000000000","0000000111000001110000011100","0000010010010100100101001001","0000011111110111111101111111","0000111000101110001011100010","0000110101011101010111010101","0000110100011101000111010001","0000101011111010111110101111","0000100110111001101110011011","0000100011001000110010001100","0000101001111010011110100111","0000101000101010001010100010","0000100110101001101010011010","0000101111101011111010111110","0000110000011100000111000001","0000101111101011111010111110","0000101111101011111010111110","0000110010101100101011001010","0000110100101101001011010010","0000100111111001111110011111","0000010001010100010101000101","0001000000000000000000000000","0001000000000000000000000000","0000000001000000010000000100","0000000100010001000100010001","0000000101100001011000010110","0000010001000100010001000100","0000100101101001011010010110","0000110011111100111111001111","0000111010101110101011101010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111100011111000111110001","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000111101101111011011110110","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111100001111000011110000","0000110010111100101111001011","0000011000010110000101100001","0000000011110000111100001111","0000000011010000110100001101","0000100010001000100010001000","0000011101000111010001110100","0000101000101010001010100010","0000011011010110110101101101","0000001011100010111000101110","0000010100110101001101010011","0000011111110111111101111111","0000100110011001100110011001","0000101101001011010010110100","0000111000001110000011100000","0000101010011010100110101001","0000110101011101010111010101","0000110111011101110111011101","0000101110011011100110111001","0000101000011010000110100001","0000011011100110111001101110","0000101111011011110110111101","0000100110011001100110011001","0000100010101000101010001010","0000011001110110011101100111","0001000000000000000000000000","0000101101101011011010110110","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000101001101010011010100110","0001000000000000000000000000","0000001111000011110000111100","0000010100000101000001010000","0000011100010111000101110001","0000100101101001011010010110","0000011100010111000101110001","0000100011011000110110001101","0000100101101001011010010110","0000100010111000101110001011","0000100101001001010010010100","0000101001101010011010100110","0000111000011110000111100001","0000111110011111100111111001","0000111111111111111111111111","0000110110011101100111011001","0000111100111111001111110011","0000110110001101100011011000","0000111100001111000011110000","0000111011111110111111101111","0000101100001011000010110000","0000100010101000101010001010","0000010100110101001101010011","0000010011110100111101001111","0000100000011000000110000001","0000101001111010011110100111","0000101000011010000110100001","0000011100000111000001110000","0000001001000010010000100100","0001000000000000000000000000","0000000010010000100100001001","0000100110001001100010011000","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111110101111101011111010","0000111110111111101111111011","0000111010101110101011101010","0000110100101101001011010010","0000101000011010000110100001","0000010001110100011101000111","0001000000000000000000000000","0001000000000000000000000000","0000000000010000000100000001","0000001110110011101100111011","0000000111010001110100011101","0000011101000111010001110100","0000011000110110001101100011","0000011011010110110101101101","0000010000110100001101000011","0000011100110111001101110011","0000111011001110110011101100","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000101001101010011010100110","0000101110011011100110111001","0000011011100110111001101110","0000110110101101101011011010","0000100101001001010010010100","0000100011001000110010001100","0000001100110011001100110011","0000001000010010000100100001","0000111000111110001111100011","0000111111111111111111111111","0000111110011111100111111001","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000101110101011101010111010","0000000001000000010000000100","0000001100010011000100110001","0000001011110010111100101111","0000001010000010100000101000","0000011100010111000101110001","0000100101111001011110010111","0000100000001000000010000000","0000100111111001111110011111","0000101101101011011010110110","0000101111101011111010111110","0000101111001011110010111100","0000100011111000111110001111","0000100011111000111110001111","0000101100111011001110110011","0000111011101110111011101110","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111110011111100111111001","0000110010011100100111001001","0000011100010111000101110001","0000001100010011000100110001","0000011110000111100001111000","0000101101101011011010110110","0000100111101001111010011110","0000110001111100011111000111","0000111110001111100011111000","0000111111001111110011111100","0000111111001111110011111100","0000110010001100100011001000","0000011000000110000001100000","0001000000000000000000000000","0000000100100001001000010010","0000010100100101001001010010","0000010111000101110001011100","0000011001000110010001100100","0000101001001010010010100100","0000110101111101011111010111","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111011111110111111101111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111100111111001111110011","0000111101101111011011110110","0000111111111111111111111111","0000101110111011101110111011","0000010110110101101101011011","0000000100110001001100010011","0001000000000000000000000000","0001000000000000000000000000","0000000000100000001000000010","0000000011000000110000001100","0001000000000000000000000000","0000010100000101000001010000","0000001110100011101000111010","0000000110000001100000011000","0000001000010010000100100001","0000010011010100110101001101","0000001011110010111100101111","0000011000000110000001100000","0000100110101001101010011010","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111011101110111011101110","0000111111001111110011111100","0000111101111111011111110111","0000111101011111010111110101","0000101001101010011010100110","0000101011101010111010101110","0000010111100101111001011110","0000100010001000100010001000","0000110010101100101011001010","0000100010001000100010001000","0001000000000000000000000000","0000011010100110101001101010","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111000101110001011100010","0000000100000001000000010000","0000001001010010010100100101","0000010110000101100001011000","0000001001110010011100100111","0000001110100011101000111010","0000010100100101001001010010","0000100000011000000110000001","0000111100101111001011110010","0000100101011001010110010101","0000110100111101001111010011","0000110110111101101111011011","0000101000101010001010100010","0000010010010100100101001001","0000010000000100000001000000","0000010011110100111101001111","0000011010000110100001101000","0000101001011010010110100101","0000101100001011000010110000","0000111100011111000111110001","0000101010001010100010101000","0000010101000101010001010100","0000010010000100100001001000","0000010110000101100001011000","0000110100011101000111010001","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111011101110111011101110","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000011110100111101001111010","0000010010110100101101001011","0001000000000000000000000000","0001000000000000000000000000","0000011001000110010001100100","0000011011000110110001101100","0000000001100000011000000110","0000000010100000101000001010","0000101100001011000010110000","0000110111101101111011011110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000110110011101100111011001","0000100000011000000110000001","0000001110000011100000111000","0001000000000000000000000000","0001000000000000000000000000","0000000011100000111000001110","0000010000110100001101000011","0000010111010101110101011101","0000010100000101000001010000","0000010001010100010101000101","0000010010110100101101001011","0000011010010110100101101001","0001000000000000000000000000","0001000000000000000000000000","0000001011100010111000101110","0000010010100100101001001010","0000010001010100010101000101","0000010011100100111001001110","0000011110100111101001111010","0000101100111011001110110011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000110101001101010011010100","0000100010001000100010001000","0000100000111000001110000011","0000101000011010000110100001","0000100000101000001010000010","0000111000011110000111100001","0000010111100101111001011110","0000000001000000010000000100","0000110011101100111011001110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000100001001000010010000100","0000000110000001100000011000","0000010001010100010101000101","0000011011000110110001101100","0000011111100111111001111110","0000110010111100101111001011","0000010001110100011101000111","0000011000010110000101100001","0000001110010011100100111001","0000100010011000100110001001","0000100111101001111010011110","0000101000111010001110100011","0000101000011010000110100001","0000011101000111010001110100","0000010110100101101001011010","0000001111100011111000111110","0000001111000011110000111100","0000000000100000001000000010","0000000000010000000100000001","0001000000000000000000000000","0000010100010101000101010001","0000010100100101001001010010","0000001111010011110100111101","0000110000011100000111000001","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111010001110100011101000","0000110010111100101111001011","0000110010011100100111001001","0000100101101001011010010110","0000001100010011000100110001","0000001111010011110100111101","0000011000000110000001100000","0000000000110000001100000011","0000000100010001000100010001","0000100011101000111010001110","0000100001101000011010000110","0001000000000000000000000000","0000010110000101100001011000","0000110001111100011111000111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111100011111000111110001","0000111011111110111111101111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111110001111100011111000","0000111110111111101111111011","0000111110101111101011111010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110010001100100011001000","0000010110100101101001011010","0000000001010000010100000101","0001000000000000000000000000","0000011100100111001001110010","0000100110001001100010011000","0000101010101010101010101010","0000110100011101000111010001","0000110101111101011111010111","0000111000101110001011100010","0000110011011100110111001101","0000110100001101000011010000","0000110010101100101011001010","0000000010100000101000001010","0000010101110101011101010111","0000011000110110001101100011","0000010110010101100101011001","0000011100110111001101110011","0000001101010011010100110101","0000010110100101101001011010","0000011110000111100001111000","0000100010011000100110001001","0000111100111111001111110011","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000101110101011101010111010","0000010001000100010001000100","0000001011010010110100101101","0000100001111000011110000111","0000101101001011010010110100","0000101100001011000010110000","0000000100000001000000010000","0000011010000110100001101000","0000111111111111111111111111","0000111110101111101011111010","0000111100101111001011110010","0000111010101110101011101010","0000000001000000010000000100","0000001110010011100100111001","0000010110000101100001011000","0000101101001011010010110100","0000110110101101101011011010","0000111101001111010011110100","0000011101100111011001110110","0000010101110101011101010111","0000001000010010000100100001","0000010001000100010001000100","0000110111101101111011011110","0000111101111111011111110111","0000101111011011110110111101","0000100001011000010110000101","0000100100011001000110010001","0000101000011010000110100001","0000100010111000101110001011","0000011000110110001101100011","0000011101110111011101110111","0000010111100101111001011110","0000001010100010101000101010","0000000001000000010000000100","0000011101110111011101110111","0000110011011100110111001101","0000111111111111111111111111","0000111001011110010111100101","0000111011011110110111101101","0000111011011110110111101101","0000111011001110110011101100","0000111101101111011011110110","0000111100011111000111110001","0000101111001011110010111100","0000011111100111111001111110","0000000110100001101000011010","0000010101000101010001010100","0000100000101000001010000010","0000101001011010010110100101","0000101110001011100010111000","0000011010000110100001101000","0000010001000100010001000100","0000101110111011101110111011","0000101001101010011010100110","0000001101000011010000110100","0000000110010001100100011001","0000110111101101111011011110","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111100011111000111110001","0000111111101111111011111110","0000111111111111111111111111","0000111101111111011111110111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111110011111100111111001","0000111111011111110111111101","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110001101100011011000","0000100111011001110110011101","0000010101000101010001010100","0000000100100001001000010010","0000010100010101000101010001","0000101011001010110010101100","0000110111101101111011011110","0000111011111110111111101111","0000111010111110101111101011","0000110111101101111011011110","0000101101101011011010110110","0000100101101001011010010110","0000100101101001011010010110","0000100111101001111010011110","0000011101010111010101110101","0000001111110011111100111111","0000010110100101101001011010","0000010001100100011001000110","0000011000100110001001100010","0000100000111000001110000011","0000001011100010111000101110","0000101010001010100010101000","0000110110001101100011011000","0000010110100101101001011010","0000010101110101011101010111","0000101100101011001010110010","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111101111111011111110111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111001011110010111100101","0000010110000101100001011000","0000000011010000110100001101","0000011100110111001101110011","0000100100101001001010010010","0000101001011010010110100101","0000010010000100100001001000","0000000010000000100000001000","0000111010001110100011101000","0000111111011111110111111101","0000111111111111111111111111","0000011010010110100101101001","0000000101000001010000010100","0000001100100011001000110010","0000100001011000010110000101","0000110100011101000111010001","0000111100001111000011110000","0000111111111111111111111111","0000101011111010111110101111","0000010110000101100001011000","0000010001010100010101000101","0000000110110001101100011011","0000011110000111100001111000","0000110001011100010111000101","0000100111011001110110011101","0000100111111001111110011111","0000100000011000000110000001","0000100000111000001110000011","0000100100101001001010010010","0000101011001010110010101100","0000100000011000000110000001","0000011010110110101101101011","0000000011000000110000001100","0000011101100111011001110110","0000100100001001000010010000","0000110110011101100111011001","0000111011101110111011101110","0000111010001110100011101000","0000111001111110011111100111","0000111011101110111011101110","0000111001011110010111100101","0000100111001001110010011100","0000001101110011011100110111","0000001011010010110100101101","0000011100100111001001110010","0000110000001100000011000000","0000100100111001001110010011","0000011111110111111101111111","0000011011000110110001101100","0000011000010110000101100001","0000011010110110101101101011","0000010101110101011101010111","0000100010101000101010001010","0000110111111101111111011111","0000101011001010110010101100","0000001111100011111000111110","0000001010000010100000101000","0000111010101110101011101010","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111011011110110111101101","0000111101101111011011110110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111110011111100111111001","0000111001011110010111100101","0000110000001100000011000000","0000011101100111011001110110","0001000000000000000000000000","0000000001010000010100000101","0000011001010110010101100101","0000100010001000100010001000","0000101011011010110110101101","0000101000111010001110100011","0000110001001100010011000100","0000110001101100011011000110","0000101011111010111110101111","0000111011101110111011101110","0000110010011100100111001001","0000101100001011000010110000","0000101110111011101110111011","0000101100011011000110110001","0000011001100110011001100110","0000011000000110000001100000","0000100001001000010010000100","0000011101000111010001110100","0000010111100101111001011110","0000011110100111101001111010","0000101110111011101110111011","0000111001111110011111100111","0000101101101011011010110110","0000100010101000101010001010","0000010010010100100101001001","0000011010000110100001101000","0000111101011111010111110101","0000111011011110110111101101","0000111011011110110111101101","0000111101101111011011110110","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000100001001000010010000100","0000000011100000111000001110","0000011010010110100101101001","0000011101010111010101110101","0000100001111000011110000111","0000101011011010110110101101","0001000000000000000000000000","0000101110101011101010111010","0000111111111111111111111111","0000111010111110101111101011","0000001010100010101000101010","0000001011000010110000101100","0000011011000110110001101100","0000101100101011001010110010","0000111010011110100111101001","0000111111011111110111111101","0000111111111111111111111111","0000111010101110101011101010","0000011100110111001101110011","0000010010010100100101001001","0000001111000011110000111100","0000001100000011000000110000","0000001111010011110100111101","0000100011011000110110001101","0000011011100110111001101110","0000011010110110101101101011","0000011110100111101001111010","0000011111100111111001111110","0000010101010101010101010101","0000001011000010110000101100","0000001001100010011000100110","0000100011101000111010001110","0000110000101100001011000010","0000110010101100101011001010","0000111100101111001011110010","0000110001011100010111000101","0000101101101011011010110110","0000101011111010111110101111","0000011101110111011101110111","0000010010000100100001001000","0000011010100110101001101010","0000101100111011001110110011","0000111000001110000011100000","0000111011111110111111101111","0000110101111101011111010111","0000101101111011011110110111","0000101000111010001110100011","0000011010000110100001101000","0000011000000110000001100000","0000010110000101100001011000","0000011001000110010001100100","0000011001000110010001100100","0000100000101000001010000010","0000111111111111111111111111","0000101001011010010110100101","0000000000010000000100000001","0000011011100110111001101110","0000111100011111000111110001","0000111111111111111111111111","0000111100101111001011110010","0000111011101110111011101110","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111110001111100011111000","0000111011011110110111101101","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111101001111010011110100","0000111110101111101011111010","0000111101101111011011110110","0000111101101111011011110110","0000111110111111101111111011","0000111010001110100011101000","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000100110111001101110011011","0000001010000010100000101000","0001000000000000000000000000","0001000000000000000000000000","0000001101000011010000110100","0000010111010101110101011101","0000010011000100110001001100","0000001011110010111100101111","0000010010100100101001001010","0000100111101001111010011110","0000101001101010011010100110","0000100011111000111110001111","0000111011011110110111101101","0000111001001110010011100100","0000110110111101101111011011","0000111001111110011111100111","0000110101101101011011010110","0000110000011100000111000001","0000100110011001100110011001","0000100001111000011110000111","0000101011111010111110101111","0000101000101010001010100010","0000101011101010111010101110","0000101010111010101110101011","0000111101111111011111110111","0000111101101111011011110110","0000111000011110000111100001","0000100101011001010110010101","0000010100110101001101010011","0000010010010100100101001001","0000100110101001101010011010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111010101110101011101010","0000111111011111110111111101","0000101011011010110110101101","0000001000110010001100100011","0000010110110101101101011011","0000011101010111010101110101","0000100001101000011010000110","0000100110011001100110011001","0000010110010101100101011001","0000011010010110100101101001","0000111110101111101011111010","0000110100011101000111010001","0000000001000000010000000100","0000011000010110000101100001","0000101100011011000110110001","0000101111111011111110111111","0000111011011110110111101101","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000101101011011010110110101","0000011010000110100001101000","0000010011010100110101001101","0000001101000011010000110100","0000010011010100110101001101","0000000011110000111100001111","0001000000000000000000000000","0000000011010000110100001101","0001000000000000000000000000","0000000100110001001100010011","0000000110000001100000011000","0000010100110101001101010011","0000101000011010000110100001","0000101000011010000110100001","0000110110111101101111011011","0000111011001110110011101100","0000101010011010100110101001","0000011110100111101001111010","0000010101000101010001010100","0000001110110011101100111011","0000010110000101100001011000","0000101011111010111110101111","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111110101111101011111010","0000111011101110111011101110","0000011010100110101001101010","0000001111110011111100111111","0000011110000111100001111000","0000010011100100111001001110","0000001100000011000000110000","0000001110010011100100111001","0000011001110110011101100111","0000011001010110010101100101","0000100011111000111110001111","0000000110100001101000011010","0000000001010000010100000101","0000001111000011110000111100","0000100010011000100110001001","0000110010001100100011001000","0000111111011111110111111101","0000111100011111000111110001","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000100001101000011010000110","0000000010010000100100001001","0001000000000000000000000000","0000010110100101101001011010","0000011001110110011101100111","0000001001100010011000100110","0000001111000011110000111100","0000010101110101011101010111","0000001011110010111100101111","0000000011000000110000001100","0000001101010011010100110101","0000010001000100010001000100","0000011111010111110101111101","0000111000111110001111100011","0000011111110111111101111111","0000011110110111101101111011","0000011111110111111101111111","0000100111001001110010011100","0000110101001101010011010100","0000110001101100011011000110","0000110000011100000111000001","0000110110111101101111011011","0000110110101101101011011010","0000111111111111111111111111","0000110110001101100011011000","0000110110011101100111011001","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000110110011101100111011001","0000011100100111001001110010","0000001111010011110100111101","0000000011110000111100001111","0000100011011000110110001101","0000111101011111010111110101","0000111101011111010111110101","0000111100101111001011110010","0000111100101111001011110010","0000111011101110111011101110","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000110000111100001111000011","0000001011100010111000101110","0000001100100011001000110010","0000011001100110011001100110","0000011110110111101101111011","0000011011000110110001101100","0000100101011001010110010101","0000000111000001110000011100","0000111110101111101011111010","0000100001111000011110000111","0000000100100001001000010010","0000011100100111001001110010","0000110001001100010011000100","0000110011001100110011001100","0000110111011101110111011101","0000111111111111111111111111","0000111100011111000111110001","0000111101001111010011110100","0000111100011111000111110001","0000110010011100100111001001","0000101010011010100110101001","0000011010100110101001101010","0000011110000111100001111000","0000100101011001010110010101","0000100010011000100110001001","0000100100011001000110010001","0000101110011011100110111001","0000100001011000010110000101","0000100000011000000110000001","0000100110001001100010011000","0000100101101001011010010110","0000100000111000001110000011","0000111100111111001111110011","0000110111101101111011011110","0000011110000111100001111000","0000000001110000011100000111","0000000000110000001100000011","0000001111100011111000111110","0000101101001011010010110100","0000111111101111111011111110","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000011101000111010001110100","0000001001100010011000100110","0000011111010111110101111101","0000011101110111011101110111","0000101011001010110010101100","0000101110011011100110111001","0000100100111001001110010011","0000011010110110101101101011","0000010001010100010101000101","0000001100000011000000110000","0000011000110110001101100011","0001000000000000000000000000","0001000000000000000000000000","0000000001110000011100000111","0000000011110000111100001111","0000000110010001100100011001","0000101100001011000010110000","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111001011110010111100101","0000101010001010100010101000","0000001001010010010100100101","0000000101000001010000010100","0000010110000101100001011000","0000100010001000100010001000","0000100010111000101110001011","0000011100000111000001110000","0000011101100111011001110110","0000001111000011110000111100","0001000000000000000000000000","0000001001100010011000100110","0000011100010111000101110001","0000011111110111111101111111","0000110001011100010111000101","0000111101011111010111110101","0000101000101010001010100010","0000101010111010101110101011","0000101100101011001010110010","0000111100111111001111110011","0000111111101111111011111110","0000111011011110110111101101","0000110111101101111011011110","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000110100111101001111010011","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111101111111011111110","0000111110001111100011111000","0000110110111101101111011011","0000010111110101111101011111","0000000010110000101100001011","0000011001010110010101100101","0000100101011001010110010101","0000111101001111010011110100","0000111101101111011011110110","0000111011101110111011101110","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000110110101101101011011010","0000010100010101000101010001","0000000111000001110000011100","0000001100110011001100110011","0000010101000101010001010100","0000011111000111110001111100","0000011111010111110101111101","0001000000000000000000000000","0000110111001101110011011100","0000010100100101001001010010","0000010011010100110101001101","0000010110000101100001011000","0000110011101100111011001110","0000111001101110011011100110","0000110010001100100011001000","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000110110111101101111011011","0000101101001011010010110100","0000101111011011110110111101","0000110100101101001011010010","0000101010101010101010101010","0000101010001010100010101000","0000011111110111111101111111","0000101010001010100010101000","0000100100001001000010010000","0000100000101000001010000010","0000110001101100011011000110","0000111101111111011111110111","0000111110011111100111111001","0000110001111100011111000111","0000000001100000011000000110","0000000010110000101100001011","0000010000110100001101000011","0000100000111000001110000011","0000111010111110101111101011","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111110001111100011111000","0000110010111100101111001011","0000001100000011000000110000","0000010100010101000101010001","0000101011111010111110101111","0000111000111110001111100011","0000111101011111010111110101","0000111100101111001011110010","0000111101101111011011110110","0000111011011110110111101101","0000101101111011011110110111","0000110100101101001011010010","0000011111110111111101111111","0000000010100000101000001010","0000001011110010111100101111","0000010010100100101001001010","0000000111000001110000011100","0000001001100010011000100110","0001000000000000000000000000","0001000000000000000000000000","0000100011011000110110001101","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111101111111011111110111","0000111011111110111111101111","0000111111111111111111111111","0000110001101100011011000110","0000010000100100001001000010","0001000000000000000000000000","0000001000110010001100100011","0000011101100111011001110110","0000101110011011100110111001","0000111000001110000011100000","0000111100101111001011110010","0000101010011010100110101001","0000001100010011000100110001","0000000001000000010000000100","0000000111100001111000011110","0000011110100111101001111010","0000001111110011111100111111","0000111000011110000111100001","0000101111101011111010111110","0000111111111111111111111111","0000101011001010110010101100","0000101100011011000110110001","0000111010001110100011101000","0000111111001111110011111100","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111011101110111011101110","0000111011101110111011101110","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000110010101100101011001010","0000110011101100111011001110","0000101010101010101010101010","0000011101010111010101110101","0000000000110000001100000011","0000111100011111000111110001","0000101110101011101010111010","0000101110111011101110111011","0000111010101110101011101010","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111010111110101111101011","0000100001011000010110000101","0000010010110100101101001011","0000001010010010100100101001","0000001101110011011100110111","0000011001100110011001100110","0000100001111000011110000111","0000000111000001110000011100","0000011101010111010101110101","0000010011110100111101001111","0000010101010101010101010101","0000010110010101100101011001","0000110001111100011111000111","0000110101001101010011010100","0000110100101101001011010010","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000111001011110010111100101","0000111011101110111011101110","0000111100001111000011110000","0000111111111111111111111111","0000101110111011101110111011","0000110101111101011111010111","0000111111111111111111111111","0000111010101110101011101010","0000110000011100000111000001","0000111101111111011111110111","0000100001101000011010000110","0000000100000001000000010000","0000010111100101111001011110","0000010101100101011001010110","0000101101001011010010110100","0000111110101111101011111010","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000101011101010111010101110","0000001010010010100100101001","0000010010010100100101001001","0000101000011010000110100001","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000110111001101110011011100","0000110011011100110111001101","0000110110111101101111011011","0000001001000010010000100100","0000000010000000100000001000","0000010000000100000001000000","0000010011110100111101001111","0000001101100011011000110110","0000010100100101001001010010","0000011010100110101001101010","0001000000000000000000000000","0000000011000000110000001100","0000110001001100010011000100","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000101000111010001110100011","0000000000100000001000000010","0000001011010010110100101101","0000100111101001111010011110","0000110000011100000111000001","0000111010011110100111101001","0000111111111111111111111111","0000111110001111100011111000","0000111001101110011011100110","0000101101111011011110110111","0000010001010100010101000101","0000000000010000000100000001","0000010100110101001101010011","0000011011010110110101101101","0000100011001000110010001100","0000100110101001101010011010","0000111100111111001111110011","0000111110011111100111111001","0000101100001011000010110000","0000110000111100001111000011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111011001110110011101100","0000111111001111110011111100","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111110011111100111111001","0000101110101011101010111010","0000110001111100011111000111","0000110010101100101011001010","0000011011110110111101101111","0000010010000100100001001000","0000110100111101001111010011","0000110101111101011111010111","0000110000101100001011000010","0000111100101111001011110010","0000111101111111011111110111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111010101110101011101010","0000100111111001111110011111","0000100011111000111110001111","0000010101010101010101010101","0000000111000001110000011100","0000010100000101000001010000","0000011100010111000101110001","0000011001110110011101100111","0000001001000010010000100100","0000000100000001000000010000","0000010111000101110001011100","0000011000100110001001100010","0000100111101001111010011110","0000100111001001110010011100","0000111100101111001011110010","0000111111111111111111111111","0000111100011111000111110001","0000111100111111001111110011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111001111110011111100","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111011001110110011101100","0000110101001101010011010100","0000110100111101001111010011","0000111011111110111111101111","0000111010111110101111101011","0000110000001100000011000000","0000111100101111001011110010","0000011110000111100001111000","0000001011110010111100101111","0000100010011000100110001001","0000010100000101000001010000","0000110001001100010011000100","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111011011110110111101101","0000110000001100000011000000","0000100100101001001010010010","0000001101010011010100110101","0000101011111010111110101111","0000111100101111001011110010","0000111101101111011011110110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000110000001100000011000000","0000101010001010100010101000","0000001101110011011100110111","0000001110010011100100111001","0000001111000011110000111100","0000010011010100110101001101","0000001111100011111000111110","0000011000110110001101100011","0000011110000111100001111000","0000100011011000110110001101","0000010000100100001001000010","0001000000000000000000000000","0000011101100111011001110110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111110001111100011111000","0000111011101110111011101110","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000011111110111111101111111","0000000001100000011000000110","0000010001010100010101000101","0000101100101011001010110010","0000110011011100110111001101","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000101001001010010010100100","0000011010110110101101101011","0000000110000001100000011000","0000000100000001000000010000","0000001110100011101000111010","0000011011000110110001101100","0000101100001011000010110000","0000111101101111011011110110","0000110000101100001011000010","0000011111010111110101111101","0000101011011010110110101101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111001111110011111100","0000111011011110110111101101","0000100110101001101010011010","0000101011001010110010101100","0000111101001111010011110100","0000011011100110111001101110","0000000100010001000100010001","0000111100011111000111110001","0000100110101001101010011010","0000100110011001100110011001","0000111011001110110011101100","0000111111101111111011111110","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111001101110011011100110","0000110110101101101011011010","0000101111001011110010111100","0000101001011010010110100101","0001000000000000000000000000","0000001011000010110000101100","0000010101000101010001010100","0000101001101010011010100110","0000000000010000000100000001","0000001010110010101100101011","0000011010100110101001101010","0000001011000010110000101100","0000010111110101111101011111","0000101001001010010010100100","0000111100101111001011110010","0000111001101110011011100110","0000111101001111010011110100","0000111011011110110111101101","0000101111111011111110111111","0000111000101110001011100010","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111101001111010011110100","0000111110111111101111111011","0000111011101110111011101110","0000110101111101011111010111","0000110001111100011111000111","0000111111111111111111111111","0000110111101101111011011110","0000101101001011010010110100","0000111111111111111111111111","0000110010111100101111001011","0000000100010001000100010001","0000010001100100011001000110","0000011101010111010101110101","0000100001011000010110000101","0000110010111100101111001011","0000111100111111001111110011","0000110100001101000011010000","0000111110001111100011111000","0000111100111111001111110011","0000111011001110110011101100","0000110001111100011111000111","0000111010011110100111101001","0000011011110110111101101111","0000100101101001011010010110","0000111100011111000111110001","0000111101001111010011110100","0000111111111111111111111111","0000111010111110101111101011","0000111110101111101011111010","0000111111001111110011111100","0000110111001101110011011100","0000011110110111101101111011","0000010011000100110001001100","0000001011010010110100101101","0000100010011000100110001001","0000100000101000001010000010","0000011101000111010001110100","0000110000101100001011000010","0000111100111111001111110011","0000110000111100001111000011","0000100111011001110110011101","0000101101101011011010110110","0000010001010100010101000101","0000010010000100100001001000","0000111000111110001111100011","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111100111111001111110011","0000100101001001010010010100","0001000000000000000000000000","0000010111000101110001011100","0000101101111011011110110111","0000101101001011010010110100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111011001110110011101100","0000111000001110000011100000","0000110000001100000011000000","0000101000011010000110100001","0000011110010111100101111001","0000010011010100110101001101","0000001100000011000000110000","0000000011010000110100001101","0000001011000010110000101100","0000101010101010101010101010","0000110100101101001011010010","0000010111110101111101011111","0000010010010100100101001001","0000111010101110101011101010","0000111101111111011111110111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111110011111100111111001","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111011001110110011101100","0000111101001111010011110100","0000111111111111111111111111","0000111011011110110111101101","0000110010011100100111001001","0000100100011001000110010001","0000101000011010000110100001","0000110001101100011011000110","0000010100000101000001010000","0000001100110011001100110011","0000110000001100000011000000","0000011101000111010001110100","0000100000101000001010000010","0000111000101110001011100010","0000111111001111110011111100","0000111011101110111011101110","0000111111111111111111111111","0000111110001111100011111000","0000111000101110001011100010","0000110110101101101011011010","0000111000011110000111100001","0000101101001011010010110100","0000011011010110110101101101","0001000000000000000000000000","0000001110110011101100111011","0000100010111000101110001011","0000000011000000110000001100","0000001110010011100100111001","0000010111010101110101011101","0000001101000011010000110100","0000001110010011100100111001","0000100011011000110110001101","0000111010101110101011101010","0000110100111101001111010011","0000111111111111111111111111","0000111100101111001011110010","0000111010011110100111101001","0000110100101101001011010010","0000101000101010001010100010","0000101000111010001110100011","0000100111101001111010011110","0000100111101001111010011110","0000101011001010110010101100","0000101110011011100110111001","0000101010101010101010101010","0000100100011001000110010001","0000010110010101100101011001","0000100100101001001010010010","0000110101101101011011010110","0000101101101011011010110110","0000101110001011100010111000","0000111111111111111111111111","0000101111011011110110111101","0000001101100011011000110110","0000001010110010101100101011","0000100100111001001110010011","0000011111100111111001111110","0000101110111011101110111011","0000111110111111101111111011","0000110000111100001111000011","0000111111111111111111111111","0000111010101110101011101010","0000110111011101110111011101","0000110111011101110111011101","0000111011111110111111101111","0000101011101010111010101110","0000101111111011111110111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000110110111101101111011011","0000100001001000010010000100","0000011011100110111001101110","0000000001010000010100000101","0000011101100111011001110110","0000101000111010001110100011","0000011110100111101001111010","0000110100001101000011010000","0000111101001111010011110100","0000101111011011110110111101","0000100110111001101110011011","0000100001101000011010000110","0000011111000111110001111100","0000001001100010011000100110","0000001011100010111000101110","0000111010101110101011101010","0000111111111111111111111111","0000111101001111010011110100","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000100111101001111010011110","0000000001010000010100000101","0000010111110101111101011111","0000011110110111101101111011","0000101110101011101010111010","0000111100101111001011110010","0000111110001111100011111000","0000111111101111111011111110","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111001101110011011100110","0000101110011011100110111001","0000101101111011011110110111","0000100100101001001010010010","0000011101100111011001110110","0000100110111001101110011011","0000010001010100010101000101","0000001001010010010100100101","0000000001100000011000000110","0000001111000011110000111100","0000010111010101110101011101","0000011010110110101101101011","0000011101010111010101110101","0000110010011100100111001001","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111010101110101011101010","0000111111111111111111111111","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000100101011001010110010101","0000011111000111110001111100","0000100111011001110110011101","0000100101001001010010010100","0000001000100010001000100010","0000100010011000100110001001","0000011010110110101101101011","0000100000001000000010000000","0000010011100100111001001110","0000011111100111111001111110","0000100010001000100010001000","0000100110111001101110011011","0000111001001110010011100100","0000111010111110101111101011","0000110011111100111111001111","0000110100001101000011010000","0000111001001110010011100100","0000101100111011001110110011","0000110110001101100011011000","0000000001010000010100000101","0000010010000100100001001000","0000010000110100001101000011","0000000100100001001000010010","0000011001010110010101100101","0000011001100110011001100110","0000010100000101000001010000","0000001110110011101100111011","0000010100110101001101010011","0000100000001000000010000000","0000101011101010111010101110","0000110011001100110011001100","0000110110101101101011011010","0000110100101101001011010010","0000100011111000111110001111","0000101010101010101010101010","0000100101011001010110010101","0000100001101000011010000110","0000100001111000011110000111","0000100010101000101010001010","0000100010001000100010001000","0000100010011000100110001001","0000100011111000111110001111","0000011001010110010101100101","0000001101000011010000110100","0000011100100111001001110010","0000011001100110011001100110","0000100011011000110110001101","0000101111001011110010111100","0000111111111111111111111111","0000111101101111011011110110","0000100110011001100110011001","0001000000000000000000000000","0000000010110000101100001011","0000001010100010101000101010","0000010000010100000101000001","0000100100011001000110010001","0000101011011010110110101101","0000111111111111111111111111","0000110001011100010111000101","0000101100101011001010110010","0000111111111111111111111111","0000111001111110011111100111","0000110000011100000111000001","0000111000101110001011100010","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111101101111011011110110","0000100101011001010110010101","0000010101000101010001010100","0000000101110001011100010111","0000011011110110111101101111","0000101100101011001010110010","0000100011111000111110001111","0000110111111101111111011111","0000111110111111101111111011","0000111010101110101011101010","0000111001101110011011100110","0000101110101011101010111010","0000111001111110011111100111","0000101000011010000110100001","0000001111110011111100111111","0000001000100010001000100010","0000111110111111101111111011","0000111111011111110111111101","0000111011011110110111101101","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111101001111010011110100","0000111111111111111111111111","0000110100001101000011010000","0001000000000000000000000000","0000100011001000110010001100","0000101000001010000010100000","0000100001101000011010000110","0000101010001010100010101000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000111111011111110111111101","0000111010111110101111101011","0000100011111000111110001111","0000010100000101000001010000","0000100000101000001010000010","0000111001001110010011100100","0000010110110101101101011011","0000010111010101110101011101","0000001011010010110100101101","0000010011110100111101001111","0000010011000100110001001100","0000000010110000101100001011","0000011011110110111101101111","0000100010001000100010001000","0000110111001101110011011100","0000111110101111101011111010","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111011101110111011101110","0000111110111111101111111011","0000111101111111011111110111","0000101100001011000010110000","0000011101000111010001110100","0000100111101001111010011110","0000100001111000011110000111","0000000001110000011100000111","0000010011000100110001001100","0000001101000011010000110100","0000011001110110011101100111","0000001011110010111100101111","0000010001010100010101000101","0000101110001011100010111000","0000111000001110000011100000","0000110000101100001011000010","0000101100111011001110110011","0000101111101011111010111110","0000101101101011011010110110","0000111001001110010011100100","0000111011101110111011101110","0000110100111101001111010011","0000111010101110101011101010","0000011011110110111101101111","0000000001000000010000000100","0000010011000100110001001100","0001000000000000000000000000","0000011110100111101001111010","0000011001110110011101100111","0000011001000110010001100100","0000001111010011110100111101","0000011010000110100001101000","0000010010000100100001001000","0000001111000011110000111100","0000001110010011100100111001","0000010100010101000101010001","0000011011010110110101101101","0000101001001010010010100100","0000011101110111011101110111","0000010100000101000001010000","0000001100100011001000110010","0000001001000010010000100100","0000000001100000011000000110","0001000000000000000000000000","0001000000000000000000000000","0000001010000010100000101000","0000010010110100101101001011","0000001100100011001000110010","0000001011110010111100101111","0000010010110100101101001011","0000001100000011000000110000","0000010001100100011001000110","0000100011101000111010001110","0000111010001110100011101000","0000111111111111111111111111","0000110111101101111011011110","0000011110000111100001111000","0000000001000000010000000100","0000001100000011000000110000","0000000101100001011000010110","0000001010110010101100101011","0000010111100101111001011110","0000011110100111101001111010","0000010001100100011001000110","0000100011001000110010001100","0000111000111110001111100011","0000111100101111001011110010","0000111001101110011011100110","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000111011111110111111101111","0000111101011111010111110101","0000100011001000110010001100","0000001111010011110100111101","0000001010110010101100101011","0000011111000111110001111100","0000101001111010011110100111","0000101010011010100110101001","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111100001111000011110000","0000111111101111111011111110","0000110010111100101111001011","0000001010000010100000101000","0000001101100011011000110110","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000000110100001101000011010","0000011101110111011101110111","0000111011011110110111101101","0000101100101011001010110010","0000101010111010101110101011","0000100110011001100110011001","0000110110011101100111011001","0000111101111111011111110111","0000111101101111011011110110","0000111100001111000011110000","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000110000111100001111000011","0000100110101001101010011010","0000011011110110111101101111","0000100001111000011110000111","0000100011001000110010001100","0000100101111001011110010111","0000010001100100011001000110","0000011010110110101101101011","0000001101110011011100110111","0000010010000100100001001000","0000000100010001000100010001","0000001100100011001000110010","0000101000001010000010100000","0000111000111110001111100011","0000111111111111111111111111","0000111010001110100011101000","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000101110111011101110111011","0000100001101000011010000110","0000100000101000001010000010","0000010001100100011001000110","0000000111110001111100011111","0000010010100100101001001010","0000010010110100101101001011","0000001101100011011000110110","0000011110010111100101111001","0000011010010110100101101001","0000110011111100111111001111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110101111101011111010","0000111001101110011011100110","0000111000111110001111100011","0000110111101101111011011110","0000111101001111010011110100","0000111110111111101111111011","0000010110110101101101011011","0000000000010000000100000001","0000010100100101001001010010","0000000000110000001100000011","0000010111100101111001011110","0000010001010100010101000101","0000010101000101010001010100","0000010000010100000101000001","0000001100010011000100110001","0000010100110101001101010011","0000010101110101011101010111","0000011010000110100001101000","0000010111110101111101011111","0000010010100100101001001010","0000000110110001101100011011","0000000100010001000100010001","0000001100100011001000110010","0000011011110110111101101111","0000101010001010100010101000","0000101110111011101110111011","0000101100111011001110110011","0000101101101011011010110110","0000110001101100011011000110","0000100101011001010110010101","0000111000101110001011100010","0000110011101100111011001110","0000100111001001110010011100","0000101110001011100010111000","0000011101010111010101110101","0000010100010101000101010001","0000100000001000000010000000","0000011111010111110101111101","0000111011011110110111101101","0000111111111111111111111111","0000110001101100011011000110","0000001111010011110100111101","0000001101010011010100110101","0000001100010011000100110001","0000010101110101011101010111","0000100000001000000010000000","0000010111010101110101011101","0000110110011101100111011001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111011111110111111101111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000110100101101001011010010","0000011011000110110001101100","0000011010100110101001101010","0001000000000000000000000000","0000100001001000010010000100","0000101010001010100010101000","0000101111101011111010111110","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111010111110101111101011","0000111111111111111111111111","0000111001111110011111100111","0000111111011111110111111101","0000111111101111111011111110","0000111010101110101011101010","0001000000000000000000000000","0000100010101000101010001010","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000100000101000001010000010","0000001111100011111000111110","0000110101111101011111010111","0000111100101111001011110010","0000110010111100101111001011","0000100100111001001110010011","0000010101010101010101010101","0000011111000111110001111100","0000100001111000011110000111","0000100010011000100110001001","0000100010001000100010001000","0000101000111010001110100011","0000110110011101100111011001","0000111101101111011011110110","0000111110001111100011111000","0000111111001111110011111100","0000101110111011101110111011","0000011100000111000001110000","0000100001011000010110000101","0000011010110110101101101011","0000010110000101100001011000","0000011100010111000101110001","0000001000000010000000100000","0000001110100011101000111010","0000001001000010010000100100","0000010100110101001101010011","0000001110100011101000111010","0000001110110011101100111011","0000101001111010011110100111","0000111000011110000111100001","0000111110011111100111111001","0000111101111111011111110111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000110100001101000011010000","0000101111011011110110111101","0000011101010111010101110101","0000001101100011011000110110","0000001001010010010100100101","0000011011000110110001101100","0000100101001001010010010100","0000011111010111110101111101","0000111000001110000011100000","0000110011111100111111001111","0000011111000111110001111100","0000111101111111011111110111","0000111010101110101011101010","0000111111111111111111111111","0000111110001111100011111000","0000111011111110111111101111","0000111011101110111011101110","0000111111111111111111111111","0000111011011110110111101101","0000111010101110101011101010","0000111111111111111111111111","0000111101101111011011110110","0000001111010011110100111101","0000000001010000010100000101","0000011111100111111001111110","0000000000100000001000000010","0000010111000101110001011100","0000010010110100101101001011","0000001101010011010100110101","0000000011000000110000001100","0000001010000010100000101000","0000011011110110111101101111","0000011001000110010001100100","0001000000000000000000000000","0001000000000000000000000000","0000001110010011100100111001","0000100011001000110010001100","0000110111101101111011011110","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111001111110011111100","0000111011101110111011101110","0000110101101101011011010110","0000110011011100110111001101","0000110001101100011011000110","0000110000011100000111000001","0000111101101111011011110110","0000110011101100111011001110","0000111001111110011111100111","0000110001011100010111000101","0000101010111010101110101011","0000101110001011100010111000","0000110000111100001111000011","0000111011011110110111101101","0000111011001110110011101100","0000101011111010111110101111","0000010101010101010101010101","0000001010110010101100101011","0000001110010011100100111001","0000011111110111111101111111","0000010000010100000101000001","0000101100011011000110110001","0000110100001101000011010000","0000111110001111100011111000","0000111111111111111111111111","0000111010101110101011101010","0000111100001111000011110000","0000111111111111111111111111","0000111101111111011111110111","0000101000001010000010100000","0000100101001001010010010100","0000010000110100001101000011","0001000000000000000000000000","0000011001110110011101100111","0000110010001100100011001000","0000111001011110010111100101","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100011101000111010001","0001000000000000000000000000","0000110001001100010011000100","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000110001101100011011000110","0000000100100001001000010010","0000011010000110100001101000","0000111011101110111011101110","0000110001001100010011000100","0000110000001100000011000000","0000100001111000011110000111","0000001111010011110100111101","0000011000000110000001100000","0000010001100100011001000110","0000001001000010010000100100","0000010011110100111101001111","0000010101100101011001010110","0000001011000010110000101100","0000011101110111011101110111","0000101111111011111110111111","0000100000011000000110000001","0000011101000111010001110100","0000100110001001100010011000","0000010010010100100101001001","0000010111100101111001011110","0000011001000110010001100100","0000011110000111100001111000","0000011110010111100101111001","0000100001011000010110000101","0000001000100010001000100010","0000001011110010111100101111","0000010001110100011101000111","0000011001010110010101100101","0000011010100110101001101010","0000111001001110010011100100","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000110100001101000011010000","0000111000001110000011100000","0000101010001010100010101000","0000001101000011010000110100","0000010010000100100001001000","0000011110010111100101111001","0000011111100111111001111110","0000100000011000000110000001","0000111010111110101111101011","0000111011101110111011101110","0000100111011001110110011101","0000110101001101010011010100","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000111011101110111011101110","0000111111111111111111111111","0000110011101100111011001110","0000001101110011011100110111","0000000100000001000000010000","0000010111110101111101011111","0000001001110010011100100111","0000001001110010011100100111","0000101001011010010110100101","0000001110100011101000111010","0000010011010100110101001101","0000111010101110101011101010","0000011111110111111101111111","0001000000000000000000000000","0000000100100001001000010010","0000110000001100000011000000","0000111011101110111011101110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000110111101101111011011110","0000111001001110010011100100","0000111000011110000111100001","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000111100101111001011110010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000110010111100101111001011","0000100011101000111010001110","0000010001100100011001000110","0000010011010100110101001101","0000101011101010111010101110","0000011011000110110001101100","0000110100011101000111010001","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101011101010111010101110","0000101110111011101110111011","0000010101100101011001010110","0000010010110100101101001011","0000000010100000101000001010","0000100110011001100110011001","0000110101011101010111010101","0000111111111111111111111111","0000111100011111000111110001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111110011111100111111001","0000111101111111011111110111","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000100110111001101110011011","0000001000110010001100100011","0000111100111111001111110011","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000011011110110111101101111","0000000011000000110000001100","0000101001001010010010100100","0000111010011110100111101001","0000101100101011001010110010","0000110110101101101011011010","0000101110001011100010111000","0000101001111010011110100111","0000110000111100001111000011","0000110010011100100111001001","0000101100011011000110110001","0000101101001011010010110100","0000101111101011111010111110","0000100100011001000110010001","0000010010010100100101001001","0000001110010011100100111001","0000010110010101100101011001","0000011101010111010101110101","0000011111000111110001111100","0000101000111010001110100011","0000100101101001011010010110","0000100001111000011110000111","0000101101011011010110110101","0000101001111010011110100111","0000101101001011010010110100","0000010100110101001101010011","0000010010010100100101001001","0000010011010100110101001101","0000010010010100100101001001","0000011100100111001001110010","0000110110111101101111011011","0000111111111111111111111111","0000111100101111001011110010","0000111001101110011011100110","0000111111111111111111111111","0000110100101101001011010010","0000100001101000011010000110","0000100100011001000110010001","0000101101101011011010110110","0000011101110111011101110111","0000100011101000111010001110","0000101110111011101110111011","0000111110001111100011111000","0000111111111111111111111111","0000110001111100011111000111","0000101010011010100110101001","0000111110001111100011111000","0000111110101111101011111010","0000111100101111001011110010","0000111111101111111011111110","0000111110001111100011111000","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111010001110100011101000","0000101110001011100010111000","0001000000000000000000000000","0000001100100011001000110010","0000001001000010010000100100","0000000010000000100000001000","0000010001110100011101000111","0000100000111000001110000011","0000100010101000101010001010","0000101001001010010010100100","0000011001010110010101100101","0000000011010000110100001101","0000010011100100111001001110","0000101101111011011110110111","0000111101101111011011110110","0000111111111111111111111111","0000111100011111000111110001","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110001111100011111000","0000111101011111010111110101","0000110101011101010111010101","0000100001101000011010000110","0000011011100110111001101110","0000000110000001100000011000","0000101000101010001010100010","0000010100010101000101010001","0000110110011101100111011001","0000111101111111011111110111","0000111110111111101111111011","0000111110001111100011111000","0000111011011110110111101101","0000111010101110101011101010","0000110010011100100111001001","0000110100101101001011010010","0000100010111000101110001011","0000001101000011010000110100","0000001111010011110100111101","0000010100010101000101010001","0000101111111011111110111111","0000111000001110000011100000","0000111101101111011011110110","0000111110111111101111111011","0000111101101111011011110110","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111100011111000111110001","0000001100010011000100110001","0000101000101010001010100010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111011111110111111101111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000110010101100101011001010","0001000000000000000000000000","0000011111110111111101111111","0000111000111110001111100011","0000101100101011001010110010","0000111101011111010111110101","0000111101101111011011110110","0000110101101101011011010110","0000110010101100101011001010","0000101011111010111110101111","0000111000101110001011100010","0000110111001101110011011100","0000111000001110000011100000","0000101100111011001110110011","0000101100011011000110110001","0000110000101100001011000010","0000001101010011010100110101","0000011100010111000101110001","0000101000101010001010100010","0000110000011100000111000001","0000110111101101111011011110","0000111010101110101011101010","0000111100001111000011110000","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000110101011101010111010101","0000101100001011000010110000","0000011000010110000101100001","0000011001010110010101100101","0000100010001000100010001000","0000101101001011010010110100","0000111111111111111111111111","0000111011111110111111101111","0000111000001110000011100000","0000101101111011011110110111","0000101100001011000010110000","0000110100111101001111010011","0000111111101111111011111110","0000110011011100110111001101","0000101111001011110010111100","0000110110001101100011011000","0000111111001111110011111100","0000111111111111111111111111","0000111010001110100011101000","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000101010111010101110101011","0000011100010111000101110001","0000000010100000101000001010","0000001100100011001000110010","0000000111000001110000011100","0000000100110001001100010011","0000001001110010011100100111","0000011010010110100101101001","0000011010110110101101101011","0000000110100001101000011010","0000001110110011101100111011","0000100111011001110110011101","0000101010011010100110101001","0000111100111111001111110011","0000111111111111111111111111","0000111100011111000111110001","0000111100101111001011110010","0000111111101111111011111110","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111100111111001111110011","0000111110001111100011111000","0000111110011111100111111001","0000011101100111011001110110","0000010111010101110101011101","0000010110000101100001011000","0000011011010110110101101101","0000010001000100010001000100","0000100010011000100110001001","0000111000111110001111100011","0000111101011111010111110101","0000111101111111011111110111","0000111111111111111111111111","0000110111011101110111011101","0000110110011101100111011001","0000011010000110100001101000","0000000100010001000100010001","0000000110110001101100011011","0000001110010011100100111001","0000101010101010101010101010","0000101111111011111110111111","0000110101101101011011010110","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111001011110010111100101","0000100110001001100010011000","0000000100000001000000010000","0000111100001111000011110000","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000001001010010010100100101","0000001100110011001100110011","0000100101011001010110010101","0000101110001011100010111000","0000110011001100110011001100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110011011100110111001101","0000110111111101111111011111","0000101100001011000010110000","0000111010001110100011101000","0000110011101100111011001110","0000011100100111001001110010","0000111111101111111011111110","0000001010000010100000101000","0000110010011100100111001001","0000111100001111000011110000","0000111100101111001011110010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000110100011101000111010001","0000100101101001011010010110","0000011110100111101001111010","0000101010011010100110101001","0000101001101010011010100110","0000111110011111100111111001","0000110010001100100011001000","0000110101101101011011010110","0000111111001111110011111100","0000111010111110101111101011","0000110010111100101111001011","0000110000001100000011000000","0000111100001111000011110000","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111101011111010111110101","0000111001111110011111100111","0000111011101110111011101110","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111101001111010011110100","0000111111111111111111111111","0000111000011110000111100001","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000110110101101101011011010","0000100111001001110010011100","0000001010010010100100101001","0000010011010100110101001101","0000001100010011000100110001","0000001111000011110000111100","0000000001100000011000000110","0000000100010001000100010001","0000011100110111001101110011","0001000000000000000000000000","0000000101000001010000010100","0000101101011011010110110101","0000011111000111110001111100","0000111011111110111111101111","0000111111111111111111111111","0000111000111110001111100011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111110011111100111111001","0000111101001111010011110100","0000111010111110101111101011","0000111011001110110011101100","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111010111110101111101011","0000111010001110100011101000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000101000101010001010100010","0000001100000011000000110000","0000010010100100101001001010","0000100101001001010010010100","0000010111000101110001011100","0000011000000110000001100000","0000001101110011011100110111","0000101011011010110110101101","0000101111011011110110111101","0000100101011001010110010101","0000010111010101110101011101","0000000100000001000000010000","0000010010110100101101001011","0000001111010011110100111101","0000011010110110101101101011","0000100101011001010110010101","0000100100001001000010010000","0000100100001001000010010000","0000101000011010000110100001","0000110110001101100011011000","0000110011001100110011001100","0000110110111101101111011011","0000111010001110100011101000","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000100110001001100010011000","0000001101010011010100110101","0000101010111010101110101011","0000111111111111111111111111","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111100001111000011110000","0000111111111111111111111111","0000111100101111001011110010","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000100001111000011110000111","0001000000000000000000000000","0000010100000101000001010000","0000101001001010010010100100","0000100110011001100110011001","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000100000111000001110000011","0000110010001100100011001000","0000101010111010101110101011","0000101001101010011010100110","0000111110011111100111111001","0000111111011111110111111101","0000111010001110100011101000","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111101101111011011110110","0000111101011111010111110101","0000111100011111000111110001","0000111110101111101011111010","0000110011111100111111001111","0000100100111001001110010011","0000011111000111110001111100","0000101011011010110110101101","0000101101001011010010110100","0000111111111111111111111111","0000111001101110011011100110","0000111111111111111111111111","0000111001001110010011100100","0000110011011100110111001101","0000111000111110001111100011","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111101001111010011110100","0000111001101110011011100110","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111011011110110111101101","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111100111111001111110011","0000100110001001100010011000","0000010100110101001101010011","0001000000000000000000000000","0000011011100110111001101110","0000001110000011100000111000","0000001011010010110100101101","0000000100010001000100010001","0000001110100011101000111010","0000010111000101110001011100","0000000000110000001100000011","0000100001101000011010000110","0000011110010111100101111001","0000101111101011111010111110","0000111111001111110011111100","0000111010001110100011101000","0000111110111111101111111011","0000111111111111111111111111","0000111101001111010011110100","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111110011111100111111001","0000110111101101111011011110","0000110001101100011011000110","0000110001001100010011000100","0000110011011100110111001101","0000101101011011010110110101","0000111100111111001111110011","0000111111111111111111111111","0000110111111101111111011111","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111000111110001111100011","0000010110110101101101011011","0000001101100011011000110110","0000100010101000101010001010","0000010110010101100101011001","0000100101101001011010010110","0000100110011001100110011001","0000010110010101100101011001","0001000000000000000000000000","0000000001010000010100000101","0000010001110100011101000111","0000001001110010011100100111","0000000101010001010100010101","0000010101110101011101010111","0000010111010101110101011101","0000100110011001100110011001","0000100011101000111010001110","0000010010000100100001001000","0000010011110100111101001111","0000011111000111110001111100","0000101111001011110010111100","0000110001011100010111000101","0000110010001100100011001000","0000111100101111001011110010","0000110111001101110011011100","0000110111001101110011011100","0000110110011101100111011001","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000110111111101111111011111","0000010010100100101001001010","0001000000000000000000000000","0000110100111101001111010011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000110000101100001011000010","0000000010010000100100001001","0000000100110001001100010011","0000010101010101010101010101","0000100110001001100010011000","0000101010101010101010101010","0000111111111111111111111111","0000111100111111001111110011","0000111101001111010011110100","0000111111111111111111111111","0000110111101101111011011110","0000111010101110101011101010","0000111111111111111111111111","0000110100101101001011010010","0000101100001011000010110000","0000111000001110000011100000","0000011010100110101001101010","0000111111111111111111111111","0000111000001110000011100000","0000110000011100000111000001","0000110101101101011011010110","0000111010011110100111101001","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111110001111100011111000","0000111111011111110111111101","0000111111001111110011111100","0000111000111110001111100011","0000100011111000111110001111","0000100111101001111010011110","0000101010011010100110101001","0000110100101101001011010010","0000111111111111111111111111","0000111110101111101011111010","0000110110111101101111011011","0000110110111101101111011011","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111000101110001011100010","0000111110101111101011111010","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111011001110110011101100","0000110110011101100111011001","0000111111111111111111111111","0000111100001111000011110000","0000111011001110110011101100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000101011111010111110101111","0000100011001000110010001100","0001000000000000000000000000","0000000101010001010100010101","0000010101000101010001010100","0000001001110010011100100111","0000000110100001101000011010","0000000001010000010100000101","0000000110100001101000011010","0000000100010001000100010001","0000000101000001010000010100","0000100111001001110010011100","0000100101011001010110010101","0000111110101111101011111010","0000111011111110111111101111","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000110111111101111111011111","0000110110001101100011011000","0000110100101101001011010010","0000110100101101001011010010","0000110011101100111011001110","0000110000001100000011000000","0000101010111010101110101011","0000100111011001110110011101","0000100110101001101010011010","0000100100001001000010010000","0000111000101110001011100010","0000111100001111000011110000","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111101001111010011110100","0000111110111111101111111011","0000111110101111101011111010","0000001100100011001000110010","0000001101110011011100110111","0000101011011010110110101101","0000010100110101001101010011","0000101000101010001010100010","0000100000001000000010000000","0000110100111101001111010011","0000110101011101010111010101","0000101010011010100110101001","0000011110000111100001111000","0000100011001000110010001100","0000101100101011001010110010","0000011000010110000101100001","0000011100000111000001110000","0000100101011001010110010101","0000001010110010101100101011","0000001000100010001000100010","0000010011100100111001001110","0000010101000101010001010100","0000100101111001011110010111","0000110100001101000011010000","0000110110001101100011011000","0000110001001100010011000100","0000111011101110111011101110","0000111110111111101111111011","0000110101111101011111010111","0000101100011011000110110001","0000101011001010110010101100","0000110101101101011011010110","0000111111111111111111111111","0000111111111111111111111111","0000101110001011100010111000","0000100111101001111010011110","0000000111010001110100011101","0000000110010001100100011001","0000111010011110100111101001","0000111001111110011111100111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111001101110011011100110","0000111010111110101111101011","0000001010100010101000101010","0000011100110111001101110011","0000000000010000000100000001","0000011111100111111001111110","0000100110011001100110011001","0000110101011101010111010101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000011010100110101001101010","0000101100011011000110110001","0000100101101001011010010110","0000101011101010111010101110","0000100100001001000010010000","0000101000101010001010100010","0000011100010111000101110001","0000110100111101001111010011","0000101011011010110110101101","0000110001101100011011000110","0000111110011111100111111001","0000111101111111011111110111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111011111110111111101","0000111110101111101011111010","0000101010111010101110101011","0000110101101101011011010110","0000110010101100101011001010","0000111101001111010011110100","0000111101001111010011110100","0000111101101111011011110110","0000111111101111111011111110","0000111011111110111111101111","0000111111101111111011111110","0000111110101111101011111010","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000110011111100111111001111","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000110100001101000011010000","0000111110101111101011111010","0000110010001100100011001000","0000101010101010101010101010","0000011100100111001001110010","0001000000000000000000000000","0000010111010101110101011101","0000011000100110001001100010","0000001110000011100000111000","0000011000000110000001100000","0000001010000010100000101000","0000000000100000001000000010","0000010001100100011001000110","0000000111100001111000011110","0000100101111001011110010111","0000110010011100100111001001","0000110010101100101011001010","0000111010011110100111101001","0000111101001111010011110100","0000101111011011110110111101","0000011101110111011101110111","0000010101000101010001010100","0000010100010101000101010001","0000010011100100111001001110","0000001110100011101000111010","0000000101110001011100010111","0001000000000000000000000000","0000000001100000011000000110","0000001010110010101100101011","0000010011010100110101001101","0000010111110101111101011111","0000011111010111110101111101","0000100100001001000010010000","0000111111001111110011111100","0000111101001111010011110100","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000111001111110011111100111","0000001101000011010000110100","0000001000000010000000100000","0000101000001010000010100000","0000100100101001001010010010","0000011001000110010001100100","0000101000111010001110100011","0000100101011001010110010101","0000100101111001011110010111","0000110000101100001011000010","0000100111101001111010011110","0000010011110100111101001111","0000000100100001001000010010","0000000110010001100100011001","0000000011010000110100001101","0000000001000000010000000100","0000000111100001111000011110","0000001010010010100100101001","0000001100010011000100110001","0000010111010101110101011101","0000011001000110010001100100","0000100010111000101110001011","0000100011001000110010001100","0000101111001011110010111100","0000111101001111010011110100","0000111110001111100011111000","0000110111001101110011011100","0000111111111111111111111111","0000111111011111110111111101","0000110001111100011111000111","0000101011001010110010101100","0000110011011100110111001101","0000100100101001001010010010","0000100001001000010010000100","0000010001110100011101000111","0000000010100000101000001010","0000011000000110000001100000","0000111111111111111111111111","0000111100101111001011110010","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111100001111000011110000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000010101110101011101010111","0000011011000110110001101100","0000101011101010111010101110","0000010001010100010101000101","0000100100011001000110010001","0000101110111011101110111011","0000111101001111010011110100","0000111110011111100111111001","0000111111111111111111111111","0000110110001101100011011000","0000011000010110000101100001","0000011011100110111001101110","0000100100111001001110010011","0000101100001011000010110000","0000101010111010101110101011","0000010111110101111101011111","0000010011110100111101001111","0000101100001011000010110000","0000100101011001010110010101","0000101001101010011010100110","0000110111011101110111011101","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111101101111011011110110","0000111100101111001011110010","0000111100011111000111110001","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000111100001111000011110000","0000101110101011101010111010","0000110110101101101011011010","0000111001111110011111100111","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111100001111000011110000","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000110101001101010011010100","0000111110001111100011111000","0000111111111111111111111111","0000110010001100100011001000","0000111110111111101111111011","0000110010111100101111001011","0000110010001100100011001000","0000001001110010011100100111","0000010010000100100001001000","0000011000110110001101100011","0000011000010110000101100001","0000001110000011100000111000","0000010000110100001101000011","0000001010010010100100101001","0000000100110001001100010011","0000011011000110110001101100","0000010001100100011001000110","0000100010011000100110001001","0000100000011000000110000001","0000101111011011110110111101","0000111100001111000011110000","0000110001001100010011000100","0000110101001101010011010100","0000111010001110100011101000","0000111111111111111111111111","0000111011011110110111101101","0000111011011110110111101101","0000111100011111000111110001","0000111110111111101111111011","0000111110111111101111111011","0000110101101101011011010110","0000100010011000100110001001","0000010001110100011101000111","0000000101010001010100010101","0000010100010101000101010001","0000011101010111010101110101","0000101101111011011110110111","0000111110011111100111111001","0000111111111111111111111111","0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100011101000111010001","0000110001101100011011000110","0000000111100001111000011110","0000010000100100001001000010","0000010101100101011001010110","0000100011001000110010001100","0000010111000101110001011100","0000011011000110110001101100","0000010001110100011101000111","0000010010110100101101001011","0000001010000010100000101000","0000000110100001101000011010","0000001011100010111000101110","0000100011011000110110001101","0000100100101001001010010010","0000011111110111111101111111","0000010110100101101001011010","0000010100110101001101010011","0000000011100000111000001110","0000000111010001110100011101","0000001010100010101000101010","0000001101100011011000110110","0000100010111000101110001011","0000101011001010110010101100","0000100111001001110010011100","0000101100001011000010110000","0000110100001101000011010000","0000111001111110011111100111","0000111111011111110111111101","0000111010111110101111101011","0000111111111111111111111111","0000111011111110111111101111","0000111100011111000111110001","0000101100111011001110110011","0000010011000100110001001100","0000001001100010011000100110","0000000110110001101100011011","0000000011010000110100001101","0000110000111100001111000011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100101111001011110010","0000100100111001001110010011","0000001011110010111100101111","0000101110011011100110111001","0000100101111001011110010111","0000100101001001010010010100","0000011111110111111101111111","0000101111111011111110111111","0000111111111111111111111111","0000111100011111000111110001","0000110011011100110111001101","0000011000110110001101100011","0000000111100001111000011110","0000101001101010011010100110","0000101001001010010010100100","0000111111001111110011111100","0000110100101101001011010010","0000011010010110100101101001","0000010001110100011101000111","0000101010001010100010101000","0000100100011001000110010001","0000101011011010110110101101","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111010001110100011101000","0000111100001111000011110000","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000110010111100101111001011","0000110101011101010111010101","0000111101011111010111110101","0000111100011111000111110001","0000111110011111100111111001","0000111111011111110111111101","0000111011111110111111101111","0000111111111111111111111111","0000111101001111010011110100","0000111011011110110111101101","0000111011001110110011101100","0000111111111111111111111111","0000111110011111100111111001","0000111011111110111111101111","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000111101001111010011110100","0000111000011110000111100001","0000110110111101101111011011","0000110110101101101011011010","0000101111001011110010111100","0000110101101101011011010110","0000111111111111111111111111","0000111001011110010111100101","0000101001011010010110100101","0000110101111101011111010111","0000100110111001101110011011","0000001010000010100000101000","0000100001001000010010000100","0000011111010111110101111101","0000011000000110000001100000","0000001111010011110100111101","0000000001010000010100000101","0000000100000001000000010000","0000001011010010110100101101","0000010100110101001101010011","0000011101010111010101110101","0000011101010111010101110101","0000011000110110001101100011","0000101000001010000010100000","0000110110111101101111011011","0000110111011101110111011101","0000110101001101010011010100","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100001111000011110000","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111001011110010111100101","0000011011110110111101101111","0001000000000000000000000000","0000010110000101100001011000","0000100101011001010110010101","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111101101111011011110110","0000111111101111111011111110","0000111001011110010111100101","0000110010101100101011001010","0000110011001100110011001100","0000100110011001100110011001","0000010000110100001101000011","0000011100110111001101110011","0000000011000000110000001100","0000001001000010010000100100","0000010101100101011001010110","0000000111110001111100011111","0000001101000011010000110100","0000010001100100011001000110","0000010101110101011101010111","0000100001011000010110000101","0000110100111101001111010011","0000111000111110001111100011","0000110101111101011111010111","0000101001111010011110100111","0000100100111001001110010011","0000011110010111100101111001","0000001011000010110000101100","0000000011100000111000001110","0000010101010101010101010101","0000001110100011101000111010","0000001110010011100100111001","0000100111001001110010011100","0000100100111001001110010011","0000110010001100100011001000","0000101100001011000010110000","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111101011111010111110101","0000111011011110110111101101","0000111111111111111111111111","0000111000111110001111100011","0000100110011001100110011001","0000011010000110100001101000","0000000110010001100100011001","0000001011000010110000101100","0000000111000001110000011100","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000110011001100110011001100","0001000000000000000000000000","0000011101100111011001110110","0000100101101001011010010110","0000011110010111100101111001","0000100111001001110010011100","0000011000010110000101100001","0000100110111001101110011011","0000111111111111111111111111","0000111001011110010111100101","0000011000110110001101100011","0000000000110000001100000011","0000100010001000100010001000","0000100001011000010110000101","0000110000001100000011000000","0000111100101111001011110010","0000111010011110100111101001","0000011011000110110001101100","0000001010100010101000101010","0000101000101010001010100010","0000100110011001100110011001","0000110001001100010011000100","0000111110011111100111111001","0000111110011111100111111001","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111000011110000111100001","0000110011011100110111001101","0000110010001100100011001000","0000111011111110111111101111","0000111100001111000011110000","0000110111001101110011011100","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111011011110110111101101","0000110100111101001111010011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111101011111010111110101","0000111010011110100111101001","0000110101001101010011010100","0000110100111101001111010011","0000101011111010111110101111","0000101010101010101010101010","0000101110011011100110111001","0000101100001011000010110000","0000111000101110001011100010","0000101100111011001110110011","0000011110100111101001111010","0000010111010101110101011101","0000011100110111001101110011","0000011000110110001101100011","0000101010011010100110101001","0000100111111001111110011111","0000010100100101001001010010","0000001110100011101000111010","0000000110010001100100011001","0000000011010000110100001101","0000001101110011011100110111","0000011001000110010001100100","0000100011111000111110001111","0000010111110101111101011111","0000001101110011011100110111","0000100101011001010110010101","0000110000111100001111000011","0000101101011011010110110101","0000111001111110011111100111","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000011000100110001001100010","0000001011000010110000101100","0000011001010110010101100101","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000101101111011011110110111","0000101000011010000110100001","0000110111111101111111011111","0000000110110001101100011011","0000011101010111010101110101","0000011100000111000001110000","0000010001010100010101000101","0000001011100010111000101110","0000000010100000101000001010","0000001111010011110100111101","0000101000101010001010100010","0000100000101000001010000010","0000110011101100111011001110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000110111001101110011011100","0000101011001010110010101100","0000101010001010100010101000","0000011011000110110001101100","0000011011000110110001101100","0001000000000000000000000000","0000010100000101000001010000","0000100000001000000010000000","0000010111000101110001011100","0000011100100111001001110010","0000110000111100001111000011","0000011000110110001101100011","0000101000001010000010100000","0000110111011101110111011101","0000111111111111111111111111","0000111101011111010111110101","0000111110001111100011111000","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000110101101101011011010110","0000100001011000010110000101","0000010011100100111001001110","0000001011100010111000101110","0000000010110000101100001011","0000011100110111001101110011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111000111110001111100011","0000010000100100001001000010","0000001010110010101100101011","0000100101011001010110010101","0000011100100111001001110010","0000001111000011110000111100","0000011010110110101101101011","0000010110010101100101011001","0000011100110111001101110011","0000110001011100010111000101","0000011000100110001001100010","0001000000000000000000000000","0000010010010100100101001001","0000011010010110100101101001","0000011010010110100101101001","0000110111111101111111011111","0000111110101111101011111010","0000111101101111011011110110","0000011111100111111001111110","0000010000100100001001000010","0000100000011000000110000001","0000101110001011100010111000","0000110110001101100011011000","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111100011111000111110001","0000101001011010010110100101","0000101110101011101010111010","0000101110001011100010111000","0000101110011011100110111001","0000101000111010001110100011","0000110011111100111111001111","0000101111101011111010111110","0000101101101011011010110110","0000111000101110001011100010","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000101111001011110010111100","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111110101111101011111010","0000111010101110101011101010","0000101111111011111110111111","0000100111111001111110011111","0000101011101010111010101110","0000100111101001111010011110","0000011000000110000001100000","0000011100110111001101110011","0000010010100100101001001010","0000010011010100110101001101","0000010111110101111101011111","0000011011010110110101101101","0000011010100110101001101010","0000110110011101100111011001","0000101110011011100110111001","0000011111110111111101111111","0000001101000011010000110100","0000000110110001101100011011","0000000010010000100100001001","0001000000000000000000000000","0000010011000100110001001100","0000011001110110011101100111","0000100001001000010010000100","0000010110010101100101011001","0000001111000011110000111100","0000011111100111111001111110","0000011111000111110001111100","0000101000011010000110100001","0000110100101101001011010010","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111110101111101011111010","0000101010101010101010101010","0000010100010101000101010001","0000011001010110010101100101","0000111111111111111111111111","0000111011111110111111101111","0000111010111110101111101011","0000111111111111111111111111","0000110111011101110111011101","0000011110000111100001111000","0000101010111010101110101011","0000011110010111100101111001","0000000010010000100100001001","0000010111010101110101011101","0000010000110100001101000011","0000010111000101110001011100","0000010100110101001101010011","0000010000000100000001000000","0000011111000111110001111100","0000101000111010001110100011","0000111101111111011111110111","0000111111001111110011111100","0000111110001111100011111000","0000111011111110111111101111","0000111111111111111111111111","0000110100101101001011010010","0000101110111011101110111011","0000100110101001101010011010","0000100000001000000010000000","0000010111110101111101011111","0000000010100000101000001010","0000010011000100110001001100","0000101010011010100110101001","0000011111000111110001111100","0000011101100111011001110110","0000100110001001100010011000","0000011010000110100001101000","0000101011111010111110101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000110001101100011011000110","0000101001011010010110100101","0000101001011010010110100101","0000100111101001111010011110","0000011001000110010001100100","0001000000000000000000000000","0000110111101101111011011110","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111110011111100111111001","0000111111001111110011111100","0000111110001111100011111000","0000100000001000000010000000","0000010010000100100001001000","0000100001001000010010000100","0000100011101000111010001110","0000010110110101101101011011","0000000001100000011000000110","0000101000011010000110100001","0000011010010110100101101001","0000011001010110010101100101","0000001011100010111000101110","0001000000000000000000000000","0000011111010111110101111101","0000100000001000000010000000","0000010011100100111001001110","0000110101111101011111010111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000100100001001000010010000","0000000100000001000000010000","0000100100011001000110010001","0000111010011110100111101001","0000111010101110101011101010","0000101110101011101010111010","0000111011111110111111101111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111110111111101111111011","0000111110111111101111111011","0000111011011110110111101101","0000110000101100001011000010","0000011111110111111101111111","0000001110100011101000111010","0000010000010100000101000001","0000010101000101010001010100","0000010110100101101001011010","0000010111100101111001011110","0000100010111000101110001011","0000111000111110001111100011","0000111111101111111011111110","0000111011001110110011101100","0000111100001111000011110000","0000100111001001110010011100","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111011101110111011101110","0000111101111111011111110111","0000110100011101000111010001","0000100001011000010110000101","0000101000101010001010100010","0000010011000100110001001100","0000001111010011110100111101","0000001011000010110000101100","0000011000010110000101100001","0000011110110111101101111011","0000011011110110111101101111","0000100001111000011110000111","0000101111001011110010111100","0000100110001001100010011000","0000100010101000101010001010","0000000110000001100000011000","0000000010110000101100001011","0000001011010010110100101101","0000000011110000111100001111","0000010000110100001101000011","0000100001011000010110000101","0000011110100111101001111010","0000010010000100100001001000","0000001100010011000100110001","0000010111010101110101011101","0000010001110100011101000111","0000100100011001000110010001","0000110001011100010111000101","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111111101111111011111110","0000111010111110101111101011","0000010111110101111101011111","0000011101100111011001110110","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000110111001101110011011100","0000100011001000110010001100","0000011110010111100101111001","0000110000101100001011000010","0001000000000000000000000000","0000011100010111000101110001","0000011001000110010001100100","0000001001110010011100100111","0000010111100101111001011110","0000011101000111010001110100","0000101110111011101110111011","0000111010011110100111101001","0000111010011110100111101001","0000111111101111111011111110","0000111110011111100111111001","0000111111001111110011111100","0000111111011111110111111101","0000111110001111100011111000","0000111011011110110111101101","0000101011011010110110101101","0000101110101011101010111010","0000011010100110101001101010","0000010111000101110001011100","0000000100000001000000010000","0000101001011010010110100101","0000011111110111111101111111","0000010011000100110001001100","0000011000100110001001100010","0000100001111000011110000111","0000100100001001000010010000","0000110101101101011011010110","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111101111111011111110111","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000110011111100111111001111","0000101110111011101110111011","0000110000111100001111000011","0000101110001011100010111000","0000011101000111010001110100","0000011000110110001101100011","0000001101100011011000110110","0000111110111111101111111011","0000111110111111101111111011","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111011011110110111101101","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111011001110110011101100","0000111110011111100111111001","0000000000110000001100000011","0000101000001010000010100000","0000100110001001100010011000","0000010111010101110101011101","0000000110000001100000011000","0000000111110001111100011111","0000100110101001101010011010","0000011100100111001001110010","0001000000000000000000000000","0000010111010101110101011101","0000011011000110110001101100","0000100000101000001010000010","0000100111101001111010011110","0000101100101011001010110010","0000111011111110111111101111","0000111110011111100111111001","0000111111111111111111111111","0000111011101110111011101110","0000111000111110001111100011","0000000001010000010100000101","0000100001111000011110000111","0000101111011011110110111101","0000101111001011110010111100","0000101011001010110010101100","0000110111111101111111011111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100111111001111110011","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111010111110101111101011","0000110011111100111111001111","0000110010101100101011001010","0000101010001010100010101000","0000011110000111100001111000","0000011010010110100101101001","0000001111010011110100111101","0000010011010100110101001101","0000100001001000010010000100","0000100101011001010110010101","0000111100011111000111110001","0000101000111010001110100011","0000101101111011011110110111","0000110110011101100111011001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000011111110111111101111111","0000010111010101110101011101","0000011010100110101001101010","0000001110000011100000111000","0000010110100101101001011010","0000100001101000011010000110","0000101011101010111010101110","0000011111100111111001111110","0000100000011000000110000001","0000101010011010100110101001","0000011111010111110101111101","0000011110000111100001111000","0000000000100000001000000010","0000001101010011010100110101","0000001010000010100000101000","0000000100010001000100010001","0000001011000010110000101100","0000100011111000111110001111","0000100011011000110110001101","0000010001110100011101000111","0000010111110101111101011111","0000010010000100100001001000","0000010100010101000101010001","0000011000100110001001100010","0000111000011110000111100001","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111001111110011111100","0000111101101111011011110110","0000100011101000111010001110","0000100000111000001110000011","0000111111111111111111111111","0000111101011111010111110101","0000110111111101111111011111","0000101010101010101010101010","0000100100111001001110010011","0000100100111001001110010011","0001000000000000000000000000","0000100000001000000010000000","0000011011010110110101101101","0000001100000011000000110000","0000010110110101101101011011","0000011001010110010101100101","0000100111001001110010011100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000111111111111111111111111","0000100110001001100010011000","0000100000111000001110000011","0000001111100011111000111110","0000011000100110001001100010","0000011100110111001101110011","0000000101110001011100010111","0000010011110100111101001111","0000100111001001110010011100","0000011101010111010101110101","0000100101001001010010010100","0000111101101111011011110110","0000111111111111111111111111","0000111101011111010111110101","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000110100111101001111010011","0000110010001100100011001000","0000110100001101000011010000","0000110000111100001111000011","0000101001111010011110100111","0000100000011000000110000001","0000001010100010101000101010","0000010100100101001001010010","0000111111101111111011111110","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111101011111010111110101","0000100110001001100010011000","0000011001000110010001100100","0000110010011100100111001001","0000100100101001001010010010","0000011011100110111001101110","0000000111010001110100011101","0000000001110000011100000111","0000001110110011101100111011","0000000111010001110100011101","0000010000000100000001000000","0000011000110110001101100011","0000100010111000101110001011","0000100011001000110010001100","0000110001011100010111000101","0000111101101111011011110110","0000111000101110001011100010","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111101011111010111110101","0000100000101000001010000010","0000100000011000000110000001","0000101001101010011010100110","0000110011111100111111001111","0000101010001010100010101000","0000101011011010110110101101","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111010001110100011101000","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100001111000011110000","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111011111110111111101111","0000111110011111100111111001","0000111010101110101011101010","0000101000101010001010100010","0000010110010101100101011001","0000000101010001010100010101","0000100001111000011110000111","0000100101101001011010010110","0000100110011001100110011001","0000011110100111101001111010","0000100100111001001110010011","0000100111011001110110011101","0000100101101001011010010110","0000100111101001111010011110","0000001000010010000100100001","0000000100010001000100010001","0000010000000100000001000000","0000010001000100010001000100","0000011110100111101001111010","0000011101100111011001110110","0000100000111000001110000011","0000101101011011010110110101","0000011011010110110101101101","0000001110000011100000111000","0000010111000101110001011100","0001000000000000000000000000","0000001111110011111100111111","0000000010100000101000001010","0000000011100000111000001110","0000011001100110011001100110","0000011010110110101101101011","0000011100000111000001110000","0000011110100111101001111010","0000001110010011100100111001","0000010111000101110001011100","0000010000110100001101000011","0000001111110011111100111111","0000101100011011000110110001","0000111000111110001111100011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111110011111100111111001","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000110001111100011111000111","0000101110111011101110111011","0000111110101111101011111010","0000111011001110110011101100","0000110100101101001011010010","0000100110111001101110011011","0000100110101001101010011010","0001000000000000000000000000","0000100010111000101110001011","0000111000001110000011100000","0000001110000011100000111000","0000001100100011001000110010","0000010100010101000101010001","0000101101101011011010110110","0000110111001101110011011100","0000111100101111001011110010","0000111101101111011011110110","0000111100011111000111110001","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111110011111100111111001","0000111100001111000011110000","0000111111111111111111111111","0000111001111110011111100111","0000101101111011011110110111","0000011001110110011101100111","0000011101010111010101110101","0000010010110100101101001011","0000000100000001000000010000","0000000111000001110000011100","0000011011000110110001101100","0000101100111011001110110011","0000100001101000011010000110","0000110000001100000011000000","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110100011101000111010001","0000101111111011111110111111","0000101101111011011110110111","0000100110001001100010011000","0000111111111111111111111111","0000100000111000001110000011","0000010101010101010101010101","0000000001110000011100000111","0000101000111010001110100011","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111001101110011011100110","0000111100011111000111110001","0000010001100100011001000110","0000101000001010000010100000","0000110000001100000011000000","0000010110010101100101011001","0000011000100110001001100010","0000001101100011011000110110","0000001100110011001100110011","0000000110110001101100011011","0000010001000100010001000100","0000010011100100111001001110","0000010110000101100001011000","0000011110100111101001111010","0000110100011101000111010001","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000110000001100000011000000","0000110101101101011011010110","0000010000110100001101000011","0000110001111100011111000111","0000100010111000101110001011","0000101001101010011010100110","0000101100011011000110110001","0000110100011101000111010001","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111011111110111111101111","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111010111110101111101011","0000111110011111100111111001","0000111110011111100111111001","0000110010101100101011001010","0000010011110100111101001111","0000001010100010101000101010","0000001110100011101000111010","0000100011011000110110001101","0000011010000110100001101000","0000100100001001000010010000","0000011100100111001001110010","0001000000000000000000000000","0000010000010100000101000001","0000010010110100101101001011","0000010001000100010001000100","0000011010010110100101101001","0000011111110111111101111111","0000101000001010000010100000","0000110001101100011011000110","0000100111001001110010011100","0000011010110110101101101011","0000010101000101010001010100","0000001110000011100000111000","0000000001000000010000000100","0000001011110010111100101111","0000000111010001110100011101","0001000000000000000000000000","0000100001001000010010000100","0000010011010100110101001101","0000010011110100111101001111","0000010000110100001101000011","0000011011010110110101101101","0000010111110101111101011111","0000010111110101111101011111","0000001100100011001000110010","0000011111100111111001111110","0000111000011110000111100001","0000111001101110011011100110","0000111011001110110011101100","0000111101001111010011110100","0000111110111111101111111011","0000111111011111110111111101","0000111110101111101011111010","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000110011101100111011001110","0000111001111110011111100111","0000111101011111010111110101","0000110100011101000111010001","0000111001111110011111100111","0000011111100111111001111110","0000001011010010110100101101","0000100010011000100110001001","0000110110011101100111011001","0000100110001001100010011000","0000011100110111001101110011","0000010000010100000101000001","0000010001000100010001000100","0000111001111110011111100111","0000111010001110100011101000","0000110001111100011111000111","0000111111101111111011111110","0000111100011111000111110001","0000111111011111110111111101","0000111101111111011111110111","0000111101111111011111110111","0000111111011111110111111101","0000111100111111001111110011","0000111111011111110111111101","0000101110101011101010111010","0000100111001001110010011100","0000100000111000001110000011","0000010010000100100001001000","0000000000100000001000000010","0000000011010000110100001101","0000010111100101111001011110","0000101110101011101010111010","0000110100011101000111010001","0000101001001010010010100100","0000110111011101110111011101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000110101101101011011010110","0000101110111011101110111011","0000100111001001110010011100","0000100011011000110110001101","0000111111111111111111111111","0000110101001101010011010100","0000011001110110011101100111","0000010100110101001101010011","0000001001000010010000100100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111110001111100011111000","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000011000000110000001100000","0000100100011001000110010001","0000110001011100010111000101","0000100010101000101010001010","0000011001110110011101100111","0000100101101001011010010110","0000000100000001000000010000","0000010010010100100101001001","0000010010010100100101001001","0000010000100100001001000010","0000001000100010001000100010","0000101011011010110110101101","0000111000011110000111100001","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111010011110100111101001","0000111011011110110111101101","0000101110111011101110111011","0000010110010101100101011001","0000011000010110000101100001","0000101110011011100110111001","0000011110000111100001111000","0000011011010110110101101101","0000100000011000000110000001","0000110000011100000111000001","0000111111111111111111111111","0000111010011110100111101001","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111010101110101011101010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000110000001100000011000000","0000010001110100011101000111","0000010010110100101101001011","0000011000110110001101100011","0000011001010110010101100101","0001000000000000000000000000","0000100100011001000110010001","0000100011111000111110001111","0000100101011001010110010101","0000100110111001101110011011","0000101000101010001010100010","0000101100001011000010110000","0000100010011000100110001001","0000101011111010111110101111","0000101001111010011110100111","0000010001010100010101000101","0000001101100011011000110110","0000001111010011110100111101","0000000000010000000100000001","0000001010110010101100101011","0000000110110001101100011011","0001000000000000000000000000","0000010001100100011001000110","0000011010000110100001101000","0000011000010110000101100001","0000010110110101101101011011","0000010101010101010101010101","0000010110010101100101011001","0000011100100111001001110010","0000100111001001110010011100","0000000100110001001100010011","0000100101001001010010010100","0000111111111111111111111111","0000110101001101010011010100","0000111000101110001011100010","0000111101001111010011110100","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000111100101111001011110010","0000110111001101110011011100","0000111010001110100011101000","0000111010001110100011101000","0000111000011110000111100001","0000110110001101100011011000","0000011100100111001001110010","0000100000111000001110000011","0000101111011011110110111101","0000101010011010100110101001","0000110010111100101111001011","0000011100110111001101110011","0000010011110100111101001111","0000010111100101111001011110","0000100010011000100110001001","0000110001101100011011000110","0000101010001010100010101000","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111000111110001111100011","0000101001111010011110100111","0000011111110111111101111111","0000010100110101001101010011","0001000000000000000000000000","0001000000000000000000000000","0000010100100101001001010010","0000101011011010110110101101","0000111111111111111111111111","0000111010101110101011101010","0000110000111100001111000011","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111011111110111111101111","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111001011110010111100101","0000110011111100111111001111","0000101001111010011110100111","0000100101101001011010010110","0000111010111110101111101011","0000111111111111111111111111","0000101011101010111010101110","0000011110000111100001111000","0000001100000011000000110000","0000100011101000111010001110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111111001111110011111100","0000110010111100101111001011","0000000001000000010000000100","0000111011101110111011101110","0000101111111011111110111111","0000011010100110101001101010","0000100000001000000010000000","0000101010101010101010101010","0000011101000111010001110100","0000010010110100101101001011","0000010111110101111101011111","0000100000101000001010000010","0000101011101010111010101110","0000110001011100010111000101","0000111101111111011111110111","0000111111111111111111111111","0000111101001111010011110100","0000111010011110100111101001","0000111010111110101111101011","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111000111110001111100011","0000111101111111011111110111","0000111001111110011111100111","0000100001111000011110000111","0000001101010011010100110101","0000110001001100010011000100","0000101000011010000110100001","0000010110000101100001011000","0000100101001001010010010100","0000100010111000101110001011","0000111110011111100111111001","0000110010111100101111001011","0000111100111111001111110011","0000111011011110110111101101","0000110110001101100011011000","0000110001001100010011000100","0000111110011111100111111001","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111110101111101011111010","0000111100011111000111110001","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000101101111011011110110111","0000111010001110100011101000","0000010101100101011001010110","0000001010100010101000101010","0000000001010000010100000101","0000100001001000010010000100","0000100011011000110110001101","0000011111100111111001111110","0000101111101011111010111110","0000111111011111110111111101","0000110100101101001011010010","0000101100101011001010110010","0000110111001101110011011100","0000101111001011110010111100","0000010111110101111101011111","0000001111100011111000111110","0000011101000111010001110100","0000010100010101000101010001","0000000000010000000100000001","0000001001100010011000100110","0000000000010000000100000001","0000000011010000110100001101","0000001101100011011000110110","0000011101110111011101110111","0000011111110111111101111111","0000100011001000110010001100","0000010110000101100001011000","0000011011110110111101101111","0000011000100110001001100010","0000011011000110110001101100","0000010101000101010001010100","0000000110010001100100011001","0000110011011100110111001101","0000101110101011101010111010","0000110100001101000011010000","0000111010111110101111101011","0000111110111111101111111011","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111111001111110011111100","0000101111111011111110111111","0000100111011001110110011101","0000110011001100110011001100","0000100100101001001010010010","0000111100111111001111110011","0000111011111110111111101111","0000101010011010100110101001","0000001100110011001100110011","0000010010000100100001001000","0000001110000011100000111000","0000101100001011000010110000","0000101101011011010110110101","0000111111111111111111111111","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111100011111000111110001","0000110111101101111011011110","0000111110111111101111111011","0000101110111011101110111011","0000100110101001101010011010","0000010111000101110001011100","0000000100100001001000010010","0000000100000001000000010000","0000011000100110001001100010","0000101001111010011110100111","0000111111111111111111111111","0000111110011111100111111001","0000110001011100010111000101","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111011011110110111101101","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000111100001111000011110000","0000110011101100111011001110","0000011111010111110101111101","0000111111111111111111111111","0000111100001111000011110000","0000110111111101111111011111","0000011111110111111101111111","0000011010000110100001101000","0000000010110000101100001011","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111101111111011111110","0000111011101110111011101110","0000111111111111111111111111","0000010011100100111001001110","0000011110010111100101111001","0000111111111111111111111111","0000110101011101010111010101","0000100111001001110010011100","0000011101010111010101110101","0000101000101010001010100010","0000011100000111000001110000","0000100010101000101010001010","0000101001011010010110100101","0000111010001110100011101000","0000110110011101100111011001","0000111010111110101111101011","0000110110111101101111011011","0000110001111100011111000111","0000111001101110011011100110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000110000001100000011000000","0000110010111100101111001011","0000011110110111101101111011","0000001100000011000000110000","0000000011100000111000001110","0000000100100001001000010010","0000000001110000011100000111","0000011000100110001001100010","0000011110100111101001111010","0000110010011100100111001001","0000101100011011000110110001","0000111101101111011011110110","0000111111111111111111111111","0000101001001010010010100100","0000110101111101011111010111","0000111001001110010011100100","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000110111101101111011011110","0000111010011110100111101001","0000101011101010111010101110","0000110010011100100111001001","0001000000000000000000000000","0000000010000000100000001000","0000100011011000110110001101","0000010100100101001001010010","0000101011001010110010101100","0000111111111111111111111111","0000111011111110111111101111","0000111110001111100011111000","0000111010001110100011101000","0000111011001110110011101100","0000101111101011111010111110","0000110101111101011111010111","0000101011001010110010101100","0000100100001001000010010000","0000001000010010000100100001","0000000101000001010000010100","0000010000010100000101000001","0000001000010010000100100001","0000000101110001011100010111","0000010100010101000101010001","0000010010100100101001001010","0000101001101010011010100110","0000100101011001010110010101","0000101000101010001010100010","0000011111010111110101111101","0000101001111010011110100111","0000100011101000111010001110","0000100010111000101110001011","0000000110000001100000011000","0000001010110010101100101011","0000101010111010101110101011","0000110001011100010111000101","0000111001101110011011100110","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000110100101101001011010010","0000101011101010111010101110","0000101101011011010110110101","0000100011001000110010001100","0000111111111111111111111111","0000111101001111010011110100","0000111010001110100011101000","0000100111101001111010011110","0000010001100100011001000110","0000010110000101100001011000","0000001010000010100000101000","0000100011001000110010001100","0000101110111011101110111011","0000111101111111011111110111","0000111111011111110111111101","0000111100101111001011110010","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000101100011011000110110001","0000101001111010011110100111","0000011001010110010101100101","0000010001000100010001000100","0000000000110000001100000011","0000011101000111010001110100","0000101011101010111010101110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000110111001101110011011100","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111101101111011011110110","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111011111110111111101111","0000011111110111111101111111","0000111011101110111011101110","0000111111111111111111111111","0000111011001110110011101100","0000100000101000001010000010","0000001111010011110100111101","0000000111100001111000011110","0000101001111010011110100111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000101110111011101110111011","0001000000000000000000000000","0000101111101011111010111110","0000100110001001100010011000","0000011000100110001001100010","0000011010000110100001101000","0000011100000111000001110000","0000100100011001000110010001","0000101010011010100110101001","0000101100101011001010110010","0000110110101101101011011010","0000101110101011101010111010","0000111000101110001011100010","0000111010011110100111101001","0000111101111111011111110111","0000111110011111100111111001","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000101110001011100010111000","0000100101001001010010010100","0000011110010111100101111001","0000010111000101110001011100","0001000000000000000000000000","0001000000000000000000000000","0001000000000000000000000000","0000001101110011011100110111","0000010100010101000101010001","0000101001011010010110100101","0000100100101001001010010010","0000111100111111001111110011","0000101010111010101110101011","0000110011111100111111001111","0000110000111100001111000011","0000111001001110010011100100","0000111110101111101011111010","0000111111111111111111111111","0000111100001111000011110000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000101100111011001110110011","0000101110001011100010111000","0000101001011010010110100101","0000010110110101101101011011","0001000000000000000000000000","0000001111110011111100111111","0000010110010101100101011001","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000100111101001111010011110","0000101101011011010110110101","0000000111100001111000011110","0000000010110000101100001011","0000010001000100010001000100","0000000110010001100100011001","0000000111110001111100011111","0000010000110100001101000011","0000100100011001000110010001","0000101101011011010110110101","0000111111111111111111111111","0000111111111111111111111111","0000110101011101010111010101","0000111011111110111111101111","0000111011111110111111101111","0000110001011100010111000101","0000100101001001010010010100","0000000011010000110100001101","0000010011010100110101001101","0000100010111000101110001011","0000101110011011100110111001","0000111111111111111111111111","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000101000001010000010100000","0000100001111000011110000111","0000101000101010001010100010","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000110000001100000011000000","0000010001100100011001000110","0000010010010100100101001001","0000001010010010100100101001","0000011111110111111101111111","0000110100111101001111010011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111010101110101011101010","0000111110001111100011111000","0000101011001010110010101100","0000011001100110011001100110","0000011100010111000101110001","0000000111010001110100011101","0000011010010110100101101001","0000100111101001111010011110","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111110101111101011111010","0000110101111101011111010111","0000111011001110110011101100","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100101111001011110010","0000111110101111101011111010","0000111111001111110011111100","0000111110101111101011111010","0000111101111111011111110111","0000111111011111110111111101","0000111110101111101011111010","0000101101101011011010110110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000100110101001101010011010","0000001100000011000000110000","0000010000010100000101000001","0000001101000011010000110100","0000111011001110110011101100","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111011101110111011101110","0000001111100011111000111110","0001000000000000000000000000","0000001000100010001000100010","0000110001111100011111000111","0000101110001011100010111000","0000100001101000011010000110","0000111001001110010011100100","0000101001101010011010100110","0000100111111001111110011111","0000101101011011010110110101","0000111111111111111111111111","0000111110101111101011111010","0000111001001110010011100100","0000110100001101000011010000","0000111010101110101011101010","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111110011111100111111001","0000111110101111101011111010","0000110110001101100011011000","0000101000011010000110100001","0000100100111001001110010011","0000011010000110100001101000","0000001000110010001100100011","0000001111100011111000111110","0000001011100010111000101110","0000001000000010000000100000","0000101011001010110010101100","0000011101010111010101110101","0000110011011100110111001101","0000100111001001110010011100","0000110101011101010111010101","0000101100111011001110110011","0000111111111111111111111111","0000111101011111010111110101","0000111101101111011011110110","0000111100111111001111110011","0000111101111111011111110111","0000111101101111011011110110","0000111101001111010011110100","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000110101001101010011010100","0000110011011100110111001101","0000100110011001100110011001","0000001100010011000100110001","0000000101100001011000010110","0000000001100000011000000110","0000011110100111101001111010","0000111111001111110011111100","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000110110001101100011011000","0000111011001110110011101100","0000100111001001110010011100","0000101111101011111010111110","0000000100000001000000010000","0000000010010000100100001001","0000010011110100111101001111","0000001001110010011100100111","0001000000000000000000000000","0000010001010100010101000101","0000100101111001011110010111","0000110001111100011111000111","0000111011101110111011101110","0000111111111111111111111111","0000111101101111011011110110","0000111011101110111011101110","0000111100011111000111110001","0000111110011111100111111001","0000111000011110000111100001","0000011001010110010101100101","0001000000000000000000000000","0000001111110011111100111111","0000100011011000110110001101","0000110010011100100111001001","0000111110011111100111111001","0000111101011111010111110101","0000111111111111111111111111","0000111101101111011011110110","0000111011001110110011101100","0000111101101111011011110110","0000111111011111110111111101","0000111101001111010011110100","0000111000111110001111100011","0000100110101001101010011010","0000011111000111110001111100","0000100000111000001110000011","0000111111111111111111111111","0000111010111110101111101011","0000111010111110101111101011","0000110100111101001111010011","0000101001111010011110100111","0000011011010110110101101101","0000001101100011011000110110","0000010010000100100001001000","0000100100101001001010010010","0000111010001110100011101000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000110100101101001011010010","0000110101001101010011010100","0000011001000110010001100100","0000010101010101010101010101","0000000010010000100100001001","0000011011000110110001101100","0000111100011111000111110001","0000111111101111111011111110","0000111010001110100011101000","0000110110001101100011011000","0000110011101100111011001110","0000110100111101001111010011","0000101111101011111010111110","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000110100001101000011010000","0000001100110011001100110011","0000010010110100101101001011","0000000010110000101100001011","0000101111001011110010111100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111011111110111111101","0000111111011111110111111101","0000100010011000100110001001","0000000001100000011000000110","0000011011010110110101101101","0000110100011101000111010001","0000110011101100111011001110","0000110100011101000111010001","0000111111111111111111111111","0000110101111101011111010111","0000110111101101111011011110","0000101100111011001110110011","0000111110111111101111111011","0000111011111110111111101111","0000111111001111110011111100","0000111100111111001111110011","0000111111011111110111111101","0000111000111110001111100011","0000111100001111000011110000","0000111011111110111111101111","0000111110011111100111111001","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111101101111011011110110","0000111101111111011111110111","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111100001111000011110000","0000101111111011111110111111","0000100101011001010110010101","0000100100111001001110010011","0000000011010000110100001101","0000000010000000100000001000","0000011000010110000101100001","0000011001100110011001100110","0000011001100110011001100110","0000110000101100001011000010","0000101001011010010110100101","0000101001101010011010100110","0000110011011100110111001101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000110001111100011111000111","0000100011111000111110001111","0000001000000010000000100000","0000001111000011110000111100","0000000001000000010000000100","0000100100001001000010010000","0000111111111111111111111111","0000111101111111011111110111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000110001011100010111000101","0000110000101100001011000010","0000100000001000000010000000","0000101001001010010010100100","0000001110000011100000111000","0001000000000000000000000000","0000001101100011011000110110","0000010000000100000001000000","0000000101010001010100010101","0000010001110100011101000111","0000011111100111111001111110","0000110101111101011111010111","0000111011111110111111101111","0000111111101111111011111110","0000111101011111010111110101","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000110011101100111011001110","0000100011111000111110001111","0000000001000000010000000100","0000001100010011000100110001","0000011110000111100001111000","0000110011011100110111001101","0000111111101111111011111110","0000111100011111000111110001","0000111111111111111111111111","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000101100001011000010110000","0000101011011010110110101101","0000010100100101001001010010","0000100110111001101110011011","0000111101011111010111110101","0000110101111101011111010111","0000101010011010100110101001","0000100010111000101110001011","0000101111001011110010111100","0000100100101001001010010010","0000000011110000111100001111","0000010100010101000101010001","0000101111001011110010111100","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111011011110110111101101","0000111010011110100111101001","0000111101111111011111110111","0000111101011111010111110101","0000100110001001100010011000","0000100111111001111110011111","0000001000000010000000100000","0000001111010011110100111101","0000011101000111010001110100","0000111110111111101111111011","0000111101101111011011110110","0000111010011110100111101001","0000110001111100011111000111","0000100101001001010010010100","0000101101111011011110110111","0000110010111100101111001011","0000110001111100011111000111","0000110110011101100111011001","0000101110001011100010111000","0000110110011101100111011001","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111010001110100011101000","0000111100111111001111110011","0000110111111101111111011111","0000111111011111110111111101","0000111101001111010011110100","0000111101001111010011110100","0000111100011111000111110001","0000111100111111001111110011","0000010100010101000101010001","0000010111100101111001011110","0000000001010000010100000101","0000011111110111111101111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101111011011110110111101","0000000000100000001000000010","0000010010000100100001001000","0000101110101011101010111010","0000110000001100000011000000","0000110000001100000011000000","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111010111110101111101011","0000101101101011011010110110","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111011001110110011101100","0000111111101111111011111110","0000111100011111000111110001","0000111011101110111011101110","0000111111111111111111111111","0000110111011101110111011101","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111001111110011111100111","0000110001011100010111000101","0000010110010101100101011001","0000010111000101110001011100","0001000000000000000000000000","0000010001110100011101000111","0000010101100101011001010110","0000100011011000110110001101","0000011100100111001001110010","0000110000101100001011000010","0000011111110111111101111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000101111111011111110111111","0000010110000101100001011000","0000001101110011011100110111","0000000101100001011000010110","0000011111100111111001111110","0000111101101111011011110110","0000111111111111111111111111","0000111101101111011011110110","0000111101111111011111110111","0000111110001111100011111000","0000111101111111011111110111","0000110110001101100011011000","0000101101101011011010110110","0000011001100110011001100110","0000011011000110110001101100","0000010001100100011001000110","0000000011010000110100001101","0000010110110101101101011011","0000001100100011001000110010","0000001001000010010000100100","0000010001010100010101000101","0000011110010111100101111001","0000111111101111111011111110","0000111111111111111111111111","0000111011101110111011101110","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000101111101011111010111110","0000100011011000110110001101","0000001010110010101100101011","0000000100000001000000010000","0000010011100100111001001110","0000101111101011111010111110","0000111010101110101011101010","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111101001111010011110100","0000111000111110001111100011","0000110110111101101111011011","0000100010011000100110001001","0000010101100101011001010110","0000011011100110111001101110","0000110011001100110011001100","0000100100101001001010010010","0000100100111001001110010011","0000101011101010111010101110","0000100011101000111010001110","0000010101010101010101010101","0000001001110010011100100111","0000011100010111000101110001","0000111101111111011111110111","0000111111101111111011111110","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111011001110110011101100","0000111001011110010111100101","0000110101001101010011010100","0000011100010111000101110001","0000101100011011000110110001","0001000000000000000000000000","0000010100100101001001010010","0000100100111001001110010011","0000111001101110011011100110","0000111111111111111111111111","0000111100011111000111110001","0000101101001011010010110100","0000011010100110101001101010","0000011100100111001001110010","0000100101001001010010010100","0000011000100110001001100010","0000101101011011010110110101","0000101111101011111010111110","0000111110011111100111111001","0000111110111111101111111011","0000111100001111000011110000","0000111101111111011111110111","0000111011101110111011101110","0000111110101111101011111010","0000110001011100010111000101","0000101101111011011110110111","0000111011011110110111101101","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000100010101000101010001010","0000011010100110101001101010","0000001111000011110000111100","0000010001000100010001000100","0000111100101111001011110010","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111011101110111011101110","0001000000000000000000000000","0000000011010000110100001101","0000011011000110110001101100","0000110000111100001111000011","0000100010101000101010001010","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111100101111001011110010","0000110111111101111111011111","0000110000011100000111000001","0000100111111001111110011111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111100111111001111110011","0000111010111110101111101011","0000110111111101111111011111","0000111001001110010011100100","0000110101101101011011010110","0000101111111011111110111111","0000110010001100100011001000","0000111011011110110111101101","0000111011111110111111101111","0000111100101111001011110010","0000111111001111110011111100","0000111011001110110011101100","0000110111011101110111011101","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000110100001101000011010000","0000101100101011001010110010","0000011000000110000001100000","0000000100110001001100010011","0000000101110001011100010111","0000001100000011000000110000","0000010100100101001001010010","0000011001010110010101100101","0000100111011001110110011101","0000011010110110101101101011","0000110001001100010011000100","0000111100101111001011110010","0000111101011111010111110101","0000111101011111010111110101","0000111110011111100111111001","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111101101111011011110110","0000100101101001011010010110","0000001001110010011100100111","0000000000100000001000000010","0000010110110101101101011011","0000111000101110001011100010","0000111111101111111011111110","0000111110001111100011111000","0000111111001111110011111100","0000111110011111100111111001","0000111111011111110111111101","0000111101101111011011110110","0000110111001101110011011100","0000100000111000001110000011","0000010011110100111101001111","0000010010000100100001001000","0000000100000001000000010000","0000001101000011010000110100","0000000001110000011100000111","0000000111010001110100011101","0000001110010011100100111001","0000010101000101010001010100","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000110010101100101011001010","0000101100111011001110110011","0000011000110110001101100011","0000000010000000100000001000","0000010001100100011001000110","0000100100011001000110010001","0000110110111101101111011011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000110110001101100011011000","0000101010101010101010101010","0000011101000111010001110100","0000000011110000111100001111","0000010010110100101101001011","0000001100000011000000110000","0000001111010011110100111101","0000001010110010101100101011","0000010101010101010101010101","0000000110100001101000011010","0000010111010101110101011101","0000010001000100010001000100","0000101000011010000110100001","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111101111111011111110111","0000111111011111110111111101","0000111101101111011011110110","0000111011001110110011101100","0000110001101100011011000110","0000100110101001101010011010","0000011001100110011001100110","0000001001100010011000100110","0000010011110100111101001111","0000100101101001011010010110","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000110101101101011011010110","0000010010000100100001001000","0000000111100001111000011110","0000010000100100001001000010","0000011111100111111001111110","0000011000110110001101100011","0000011011010110110101101101","0000101101111011011110110111","0000111111111111111111111111","0000111101101111011011110110","0000111001011110010111100101","0000111011001110110011101100","0000100001011000010110000101","0000100110011001100110011001","0000110001011100010111000101","0000111010101110101011101010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000100101111001011110010111","0000010000110100001101000011","0000010110110101101101011011","0000000011000000110000001100","0000110011011100110111001101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000100101001001010010010100","0001000000000000000000000000","0000000111100001111000011110","0000101000001010000010100000","0000100011111000111110001111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111110111111101111111011","0000111100001111000011110000","0000110111001101110011011100","0000101010011010100110101001","0000111110111111101111111011","0000111111111111111111111111","0000101011001010110010101100","0000110100001101000011010000","0000111101011111010111110101","0000101000011010000110100001","0000101111001011110010111100","0000100100111001001110010011","0000011101110111011101110111","0000100111001001110010011100","0000100111111001111110011111","0000100001101000011010000110","0000101010001010100010101000","0000111011101110111011101110","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111011111110111111101","0000111100101111001011110010","0000111110001111100011111000","0000111111111111111111111111","0000111001111110011111100111","0000101100101011001010110010","0000011000010110000101100001","0000000101010001010100010101","0000001101000011010000110100","0001000000000000000000000000","0000001111100011111000111110","0000010101010101010101010101","0000011000100110001001100010","0000011000000110000001100000","0000101000011010000110100001","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000110110001101100011011000","0000100110011001100110011001","0000010111000101110001011100","0001000000000000000000000000","0000010101000101010001010100","0000110010011100100111001001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110001101100011011000110","0000011011010110110101101101","0000010110010101100101011001","0001000000000000000000000000","0000000001110000011100000111","0000001001000010010000100100","0000001110010011100100111001","0000010100110101001101010011","0000010000000100000001000000","0000111110101111101011111010","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101001111010011110100","0000111111111111111111111111","0000111011101110111011101110","0000110110111101101111011011","0000100001011000010110000101","0001000000000000000000000000","0000000110010001100100011001","0000010011010100110101001101","0000101001011010010110100101","0000111000101110001011100010","0000110111101101111011011110","0000100001001000010010000100","0000011001100110011001100110","0000000100110001001100010011","0000001111100011111000111110","0000010101010101010101010101","0000010000010100000101000001","0000001010010010100100101001","0000000100110001001100010011","0001000000000000000000000000","0000011001110110011101100111","0000100010001000100010001000","0000011011110110111101101111","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111110111111101111111011","0000111100011111000111110001","0000111000101110001011100010","0000111000101110001011100010","0000110001101100011011000110","0000101000111010001110100011","0000001010100010101000101010","0000010010100100101001001010","0000100010011000100110001001","0000100010111000101110001011","0000110111011101110111011101","0000111010101110101011101010","0000110100011101000111010001","0000011101010111010101110101","0000001011110010111100101111","0000001100110011001100110011","0000001101110011011100110111","0000010100000101000001010000","0000000100010001000100010001","0000001011100010111000101110","0000010101000101010001010100","0000011000110110001101100011","0000011000110110001101100011","0000010101000101010001010100","0000010111100101111001011110","0000110000101100001011000010","0000101011111010111110101111","0000111010011110100111101001","0000110010101100101011001010","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111111001111110011111100","0000111111011111110111111101","0000100011011000110110001101","0000001100000011000000110000","0000010111110101111101011111","0001000000000000000000000000","0000100110011001100110011001","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000010100100101001001010010","0001000000000000000000000000","0000010100100101001001010010","0000100101011001010110010101","0000111000111110001111100011","0000111001101110011011100110","0000111111111111111111111111","0000111110101111101011111010","0000110101111101011111010111","0000111101101111011011110110","0000111111111111111111111111","0000111110011111100111111001","0000110100001101000011010000","0000101101011011010110110101","0000100011011000110110001101","0000011010010110100101101001","0000101100011011000110110001","0000101101111011011110110111","0000001101110011011100110111","0000100101111001011110010111","0000101100101011001010110010","0000100111001001110010011100","0000100010011000100110001001","0000101101001011010010110100","0000111100001111000011110000","0000111011101110111011101110","0000110000011100000111000001","0000101010001010100010101000","0000111010111110101111101011","0000111111111111111111111111","0000111010111110101111101011","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111001011110010111100101","0000100110111001101110011011","0000011000110110001101100011","0001000000000000000000000000","0000010110110101101101011011","0000010111100101111001011110","0000000011000000110000001100","0000001101010011010100110101","0000010010100100101001001010","0000010011110100111101001111","0000011011100110111001101110","0000110011011100110111001101","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111100111111001111110011","0000111111101111111011111110","0000111111011111110111111101","0000111100101111001011110010","0000111110001111100011111000","0000101111001011110010111100","0000100111011001110110011101","0000100110111001101110011011","0000000010010000100100001001","0000011001010110010101100101","0000101100011011000110110001","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000101000011010000110100001","0000011100110111001101110011","0000000110100001101000011010","0000001111110011111100111111","0000010110000101100001011000","0000001100100011001000110010","0000011011010110110101101101","0000011101000111010001110100","0000110111101101111011011110","0000110011101100111011001110","0000111100101111001011110010","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111011111110111111101","0000111101111111011111110111","0000111101001111010011110100","0000111111111111111111111111","0000111011101110111011101110","0000111110011111100111111001","0000111101111111011111110111","0000100110001001100010011000","0001000000000000000000000000","0001000000000000000000000000","0000000001010000010100000101","0000000011100000111000001110","0001000000000000000000000000","0001000000000000000000000000","0000010011010100110101001101","0000011011000110110001101100","0000011111010111110101111101","0000010111000101110001011100","0000010110100101101001011010","0000011000110110001101100011","0000100111001001110010011100","0000001000110010001100100011","0000000000110000001100000011","0000000011000000110000001100","0000101111001011110010111100","0000111111111111111111111111","0000111101111111011111110111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110011111100111111001111","0000100010011000100110001001","0000011010010110100101101001","0000001000000010000000100000","0000010000110100001101000011","0000100101111001011110010111","0000100101111001011110010111","0000101011111010111110101111","0000100110101001101010011010","0000010101110101011101010111","0000010001100100011001000110","0000100100001001000010010000","0000101001101010011010100110","0000010011000100110001001100","0001000000000000000000000000","0000000101010001010100010101","0000010000100100001001000010","0000001111000011110000111100","0000000010110000101100001011","0000001001010010010100100101","0000010011010100110101001101","0000110110101101101011011010","0000111010001110100011101000","0000110100001101000011010000","0000100110111001101110011011","0000110010011100100111001001","0000111001111110011111100111","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111010011110100111101001","0000100001111000011110000111","0000010001010100010101000101","0000010011000100110001001100","0000000101100001011000010110","0000010100110101001101010011","0000111111001111110011111100","0000111111101111111011111110","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000011101110111011101110111","0000000110010001100100011001","0000100101001001010010010100","0000100010111000101110001011","0000111110001111100011111000","0000101100111011001110110011","0000110001101100011011000110","0000101010011010100110101001","0000110101111101011111010111","0000110000011100000111000001","0000100011111000111110001111","0000100000001000000010000000","0000011011010110110101101101","0000011010010110100101101001","0000010101010101010101010101","0000011100010111000101110001","0000011111010111110101111101","0000001101010011010100110101","0000001011000010110000101100","0000000100100001001000010010","0000011000100110001001100010","0000110110011101100111011001","0000111110111111101111111011","0000111111111111111111111111","0000111011101110111011101110","0000111101001111010011110100","0000111111101111111011111110","0000110000101100001011000010","0000110101011101010111010101","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111101001111010011110100","0000111110011111100111111001","0000111000111110001111100011","0000011111110111111101111111","0001000000000000000000000000","0000010011010100110101001101","0000100100001001000010010000","0000011000010110000101100001","0000001111110011111100111111","0000000010110000101100001011","0000001000100010001000100010","0000010110100101101001011010","0000010100100101001001010010","0000010110110101101101011011","0000110001001100010011000100","0000110100111101001111010011","0000110101001101010011010100","0000110011011100110111001101","0000110111101101111011011110","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111001111110011111100111","0000110001101100011011000110","0000100111111001111110011111","0001000000000000000000000000","0000011100110111001101110011","0000101001111010011110100111","0000111111101111111011111110","0000111111011111110111111101","0000111110011111100111111001","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111001001110010011100100","0000110000011100000111000001","0000101110011011100110111001","0001000000000000000000000000","0000000111110001111100011111","0000010001100100011001000110","0000000100110001001100010011","0000010001000100010001000100","0000011110010111100101111001","0000101100111011001110110011","0000101111101011111010111110","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000110100101101001011010010","0000101001011010010110100101","0000100110011001100110011001","0000100100001001000010010000","0000100001001000010010000100","0000110001011100010111000101","0000110010011100100111001001","0000100100101001001010010010","0000110000111100001111000011","0000110101011101010111010101","0000101010111010101110101011","0000101001111010011110100111","0000100101011001010110010101","0000011001000110010001100100","0000010011000100110001001100","0001000000000000000000000000","0000110000101100001011000010","0000111001101110011011100110","0000111100011111000111110001","0000111011011110110111101101","0000111011111110111111101111","0000111111111111111111111111","0000111111101111111011111110","0000101001011010010110100101","0000000110000001100000011000","0000000111010001110100011101","0000011101110111011101110111","0000011000000110000001100000","0000100100111001001110010011","0000010000100100001001000010","0000001111000011110000111100","0000001011000010110000101100","0000001011000010110000101100","0000001100000011000000110000","0000000010000000100000001000","0001000000000000000000000000","0000000011000000110000001100","0000001011000010110000101100","0000000001100000011000000110","0000000110010001100100011001","0000010010110100101101001011","0000010110000101100001011000","0000100101101001011010010110","0000100010011000100110001001","0000111010011110100111101001","0000110111101101111011011110","0000011000100110001001100010","0000100100001001000010010000","0000101011001010110010101100","0000111011001110110011101100","0000111011101110111011101110","0000111101101111011011110110","0000101000101010001010100010","0000010111100101111001011110","0000001101010011010100110101","0000000001110000011100000111","0000010011000100110001001100","0000000110110001101100011011","0000110100111101001111010011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111111011111110111111101","0000111111101111111011111110","0000010000110100001101000011","0000001100000011000000110000","0000011010110110101101101011","0000110100011101000111010001","0000100100111001001110010011","0000100000001000000010000000","0000011110000111100001111000","0000010101010101010101010101","0000001110000011100000111000","0000001101010011010100110101","0000000100000001000000010000","0000000111000001110000011100","0000001001010010010100100101","0000001011000010110000101100","0000001111110011111100111111","0000000110100001101000011010","0000001111010011110100111101","0000000011010000110100001101","0000011001000110010001100100","0000011110110111101101111011","0000111011011110110111101101","0000111100011111000111110001","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111010001110100011101000","0000111111111111111111111111","0000111011101110111011101110","0000110000101100001011000010","0000111110111111101111111011","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000110001101100011011000110","0000101101011011010110110101","0000010001000100010001000100","0000001000100010001000100010","0000101011111010111110101111","0000101000101010001010100010","0000011010000110100001101000","0000011010110110101101101011","0000001101010011010100110101","0000001000110010001100100011","0000001010110010101100101011","0000010000010100000101000001","0000011110010111100101111001","0000111000011110000111100001","0000111001101110011011100110","0000111011101110111011101110","0000111101011111010111110101","0000111110101111101011111010","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111100001111000011110000","0000011101010111010101110101","0000101001011010010110100101","0000000001110000011100000111","0000110000011100000111000001","0000110011011100110111001101","0000111011111110111111101111","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111011001110110011101100","0000111111111111111111111111","0000111101111111011111110111","0000100111111001111110011111","0000110111111101111111011111","0001000000000000000000000000","0000010000100100001001000010","0000011011010110110101101101","0000001010000010100000101000","0000000111100001111000011110","0000011000110110001101100011","0000010101110101011101010111","0000110100001101000011010000","0000111011001110110011101100","0000111011011110110111101101","0000111010101110101011101010","0000111111001111110011111100","0000111110101111101011111010","0000111001111110011111100111","0000111111111111111111111111","0000111010101110101011101010","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111100001111000011110000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111010101110101011101010","0000110001001100010011000100","0000110001101100011011000110","0000111000101110001011100010","0000110110001101100011011000","0000101111011011110110111101","0000101111111011111110111111","0000101011011010110110101101","0000100110001001100010011000","0000101010111010101110101011","0000100111011001110110011101","0000100011111000111110001111","0000100110111001101110011011","0000101011101010111010101110","0000011101110111011101110111","0000000001010000010100000101","0000111000011110000111100001","0000111011011110110111101101","0000110001011100010111000101","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000101100111011001110110011","0000000110110001101100011011","0000001001010010010100100101","0000011011100110111001101110","0000100100111001001110010011","0000011010010110100101101001","0000000000110000001100000011","0001000000000000000000000000","0000001101000011010000110100","0000000101010001010100010101","0000000111100001111000011110","0000001011110010111100101111","0000010100100101001001010010","0000100000101000001010000010","0000100100001001000010010000","0000010110010101100101011001","0000000100110001001100010011","0000000110100001101000011010","0000010001010100010101000101","0000010101110101011101010111","0000011100100111001001110010","0000001011100010111000101110","0000011101100111011001110110","0000011110110111101101111011","0000001110110011101100111011","0000001111110011111100111111","0000100011101000111010001110","0000101010001010100010101000","0000011111100111111001111110","0000010000010100000101000001","0000000100110001001100010011","0000000100000001000000010000","0000001111000011110000111100","0000101000001010000010100000","0001000000000000000000000000","0000101101001011010010110100","0000111111111111111111111111","0000111011011110110111101101","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111000001110000011100000","0000000000110000001100000011","0000010011010100110101001101","0000011110010111100101111001","0000100111111001111110011111","0000011010100110101001101010","0000100000011000000110000001","0000001101000011010000110100","0000010110110101101101011011","0000100111111001111110011111","0000110000111100001111000011","0000110111001101110011011100","0000111001101110011011100110","0000101111101011111010111110","0000110111101101111011011110","0000100110011001100110011001","0000101111001011110010111100","0000011101110111011101110111","0000000010000000100000001000","0000101000111010001110100011","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111010011110100111101001","0000111101011111010111110101","0000111111001111110011111100","0000111011111110111111101111","0000111111101111111011111110","0000111111101111111011111110","0000111010101110101011101010","0000100100001001000010010000","0000110000111100001111000011","0000101011101010111010101110","0000000010110000101100001011","0000101001101010011010100110","0000110110111101101111011011","0000100001101000011010000110","0000110100111101001111010011","0000101000101010001010100010","0000011001000110010001100100","0000010001010100010101000101","0000010001110100011101000111","0000010100110101001101010011","0000011101000111010001110100","0000110010111100101111001011","0000110100101101001011010010","0000110111101101111011011110","0000111010111110101111101011","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000100101101001011010010110","0000101100001011000010110000","0001000000000000000000000000","0000111111111111111111111111","0000111000011110000111100001","0000111110001111100011111000","0000111110011111100111111001","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111011111110111111101111","0000100101001001010010010100","0000000100100001001000010010","0000001001100010011000100110","0000100111101001111010011110","0000001000110010001100100011","0000001011110010111100101111","0000011010110110101101101011","0000001101000011010000110100","0000101011101010111010101110","0000111111111111111111111111","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111101111111011111110111","0000111001001110010011100100","0000110100111101001111010011","0000111101111111011111110111","0000110100111101001111010011","0000111110111111101111111011","0000111101101111011011110110","0000111111001111110011111100","0000111101101111011011110110","0000111001111110011111100111","0000111110111111101111111011","0000111000101110001011100010","0000111001101110011011100110","0000111001111110011111100111","0000111100001111000011110000","0000111110111111101111111011","0000111110001111100011111000","0000111101001111010011110100","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000110110111101101111011011","0000110011001100110011001100","0000101010011010100110101001","0000100111011001110110011101","0000100101001001010010010100","0000101010101010101010101010","0000010101000101010001010100","0000010110100101101001011010","0000110011101100111011001110","0000101101111011011110110111","0000110111011101110111011101","0000110100111101001111010011","0000111000001110000011100000","0000011100100111001001110010","0000001001000010010000100100","0000011000100110001001100010","0000010010100100101001001010","0000010010010100100101001001","0000000101010001010100010101","0000011110100111101001111010","0000101100101011001010110010","0000100010101000101010001010","0000010110100101101001011010","0000100010011000100110001001","0000101100111011001110110011","0000101111101011111010111110","0000101111101011111010111110","0000110001001100010011000100","0000110000001100000011000000","0000101101011011010110110101","0000011001110110011101100111","0000000001100000011000000110","0000010011110100111101001111","0000010100110101001101010011","0000010011000100110001001100","0000001110110011101100111011","0000010010110100101101001011","0000001111010011110100111101","0000001110110011101100111011","0000010010000100100001001000","0000001101010011010100110101","0000000100110001001100010011","0000001010000010100000101000","0000000100110001001100010011","0000010010000100100001001000","0000011000100110001001100010","0000100111101001111010011110","0000010110000101100001011000","0000011001000110010001100100","0000111110001111100011111000","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0001000000000000000000000000","0000001010010010100100101001","0000011110000111100001111000","0000011011110110111101101111","0000010000100100001001000010","0000100001001000010010000100","0000110110111101101111011011","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000101010001010100010101000","0000101010101010101010101010","0000101110101011101010111010","0000101010111010101110101011","0001000000000000000000000000","0000101101111011011110110111","0000111111111111111111111111","0000110111001101110011011100","0000111111111111111111111111","0000111001111110011111100111","0000111011101110111011101110","0000111011101110111011101110","0000111111111111111111111111","0000111011101110111011101110","0000110111011101110111011101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000110110101101101011011010","0000100100101001001010010010","0000100011101000111010001110","0000101011011010110110101101","0000000111110001111100011111","0000011011100110111001101110","0000110000011100000111000001","0000110010101100101011001010","0000101111101011111010111110","0000110100101101001011010010","0000101000011010000110100001","0000101111111011111110111111","0000100010011000100110001001","0000010110100101101001011010","0000100110011001100110011001","0000101001111010011110100111","0000110101101101011011010110","0000110010001100100011001000","0000101101011011010110110101","0000101010101010101010101010","0000101100101011001010110010","0000110010101100101011001010","0000111001111110011111100111","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000100111001001110010011100","0000101011111010111110101111","0000001000110010001100100011","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111011011110110111101101","0000111011001110110011101100","0000111011001110110011101100","0000101000101010001010100010","0000000011000000110000001100","0000001011000010110000101100","0000100110111001101110011011","0000010110110101101101011011","0000000111010001110100011101","0000011000100110001001100010","0000010011110100111101001111","0000011100000111000001110000","0000110111001101110011011100","0000111111111111111111111111","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111011011110110111101101","0000101110001011100010111000","0000110111001101110011011100","0000111100101111001011110010","0000110000001100000011000000","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111110011111100111111001","0000110101011101010111010101","0000100101001001010010010100","0000100010001000100010001000","0000101100001011000010110000","0000001001000010010000100100","0000100011111000111110001111","0000011110010111100101111001","0000110101011101010111010101","0000101010001010100010101000","0000100100001001000010010000","0000001100000011000000110000","0000011110000111100001111000","0000011101010111010101110101","0000000101100001011000010110","0000010101010101010101010101","0000101001101010011010100110","0000110111001101110011011100","0000101100111011001110110011","0000110011011100110111001101","0000111011011110110111101101","0000111110101111101011111010","0000111111011111110111111101","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111101111111011111110111","0000111001011110010111100101","0000110110011101100111011001","0000010111100101111001011110","0000000010000000100000001000","0000001000010010000100100001","0000010010110100101101001011","0000011001000110010001100100","0000001000010010000100100001","0000001100110011001100110011","0000001100100011001000110010","0000010001000100010001000100","0000000010110000101100001011","0000001111000011110000111100","0000011011100110111001101110","0000101010001010100010101000","0000100110101001101010011010","0000011000010110000101100001","0000011110000111100001111000","0000011011010110110101101101","0000001100000011000000110000","0000111010101110101011101010","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000110100101101001011010010","0001000000000000000000000000","0000010010110100101101001011","0000011001000110010001100100","0000001110100011101000111010","0000100001101000011010000110","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111100001111000011110000","0000111101111111011111110111","0000100010011000100110001001","0000100111001001110010011100","0000110101011101010111010101","0000000010000000100000001000","0000100011001000110010001100","0000111110011111100111111001","0000111111111111111111111111","0000111100001111000011110000","0000110110001101100011011000","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111010101110101011101010","0000110101011101010111010101","0000111010011110100111101001","0000111101011111010111110101","0000111111111111111111111111","0000111111011111110111111101","0000110111111101111111011111","0000100000111000001110000011","0000011100100111001001110010","0000101000101010001010100010","0000001010000010100000101000","0000001111110011111100111111","0000101111011011110110111101","0000110111011101110111011101","0000100111001001110010011100","0000111111011111110111111101","0000111100001111000011110000","0000110001001100010011000100","0000110001111100011111000111","0000110001101100011011000110","0000101011101010111010101110","0000111001101110011011100110","0000110011011100110111001101","0000110011001100110011001100","0000110101011101010111010101","0000111000111110001111100011","0000111100011111000111110001","0000111110101111101011111010","0000111111101111111011111110","0000111111011111110111111101","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000110001001100010011000100","0000010101010101010101010101","0000011101110111011101110111","0000111000111110001111100011","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111101011111010111110101","0000111111101111111011111110","0000111101111111011111110111","0000110111011101110111011101","0000101001101010011010100110","0000111001101110011011100110","0000001100000011000000110000","0000010001000100010001000100","0000100101111001011110010111","0000100000111000001110000011","0000010000100100001001000010","0000000100000001000000010000","0000011010110110101101101011","0000100001011000010110000101","0000101110111011101110111011","0000111010101110101011101010","0000111111111111111111111111","0000111110101111101011111010","0000111010011110100111101001","0000111111001111110011111100","0000100010111000101110001011","0000101110001011100010111000","0000111000011110000111100001","0000111011101110111011101110","0000101000101010001010100010","0000110000001100000011000000","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111110011111100111111001","0000110110001101100011011000","0000100101011001010110010101","0000100111101001111010011110","0000010100010101000101010001","0000011001110110011101100111","0000011100010111000101110001","0000100010101000101010001010","0000101010101010101010101010","0000100010011000100110001001","0000000100000001000000010000","0000100010101000101010001010","0000001000000010000000100000","0000100000101000001010000010","0000110010011100100111001001","0000110010111100101111001011","0000111001011110010111100101","0000111111101111111011111110","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000110011111100111111001111","0000100001111000011110000111","0000000001000000010000000100","0000010101000101010001010100","0000010100110101001101010011","0000010100100101001001010010","0000001101000011010000110100","0000010000100100001001000010","0000011111110111111101111111","0000101011011010110110101101","0000110001011100010111000101","0000110000111100001111000011","0000110001001100010011000100","0000111000101110001011100010","0000110111111101111111011111","0000011110010111100101111001","0000011011010110110101101101","0000000011000000110000001100","0000110100101101001011010010","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000101110101011101010111010","0001000000000000000000000000","0000010101010101010101010101","0000100000011000000110000001","0000101111011011110110111101","0000101110001011100010111000","0000111111111111111111111111","0000111101001111010011110100","0000111100101111001011110010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110011101100111011001110","0000100000001000000010000000","0000101010001010100010101000","0000010000010100000101000001","0000010010010100100101001001","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000110101111101011111010111","0000111101011111010111110101","0000111111111111111111111111","0000111100011111000111110001","0000111110001111100011111000","0000101100011011000110110001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000100101111001011110010111","0000010011100100111001001110","0000011101010111010101110101","0000000111110001111100011111","0000010100110101001101010011","0000101000101010001010100010","0000111000001110000011100000","0000011011010110110101101101","0000110101011101010111010101","0000111001011110010111100101","0000101101101011011010110110","0000110110011101100111011001","0000110001111100011111000111","0000101001111010011110100111","0000110001111100011111000111","0000111001101110011011100110","0000101010011010100110101001","0000111101001111010011110100","0000111101001111010011110100","0000111101011111010111110101","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000110111011101110111011101","0001000000000000000000000000","0000101011111010111110101111","0000110011111100111111001111","0000111011111110111111101111","0000111110001111100011111000","0000111110001111100011111000","0000111110111111101111111011","0000111101101111011011110110","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000100110001001100010011000","0000110001001100010011000100","0000010010000100100001001000","0000010010110100101101001011","0000011100110111001101110011","0000101010101010101010101010","0000100011001000110010001100","0001000000000000000000000000","0000010110000101100001011000","0000110110111101101111011011","0000100001101000011010000110","0000110011001100110011001100","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111010011110100111101001","0000100110101001101010011010","0000100001001000010010000100","0000100001101000011010000110","0000011010100110101001101010","0000100010011000100110001001","0000011110100111101001111010","0000100010011000100110001001","0000101100011011000110110001","0000111001101110011011100110","0000110111111101111111011111","0000110111101101111011011110","0000110011101100111011001110","0000110000011100000111000001","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000110001001100010011000100","0000011110100111101001111010","0000101001001010010010100100","0000100010001000100010001000","0000000111010001110100011101","0000011111100111111001111110","0000011001110110011101100111","0000011110000111100001111000","0000010001010100010101000101","0000100000111000001110000011","0000010000000100000001000000","0000100000101000001010000010","0000111111111111111111111111","0000111010111110101111101011","0000110011011100110111001101","0000111001111110011111100111","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111110011111100111111001","0000111110111111101111111011","0000111101001111010011110100","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001101110011011100110","0000011101100111011001110110","0001000000000000000000000000","0000011001110110011101100111","0000010111110101111101011111","0000011010100110101001101010","0000001010010010100100101001","0000100110011001100110011001","0000110111111101111111011111","0000110011001100110011001100","0000101000101010001010100010","0000111111111111111111111111","0000111110101111101011111010","0000110010111100101111001011","0000110000011100000111000001","0000011011100110111001101110","0000001100100011001000110010","0000011101010111010101110101","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111111101111111011111110","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000011100010111000101110001","0000001111010011110100111101","0000010110110101101101011011","0000100001101000011010000110","0000111011111110111111101111","0000111000111110001111100011","0000111100101111001011110010","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111000111110001111100011","0000110110111101101111011011","0000110010011100100111001001","0000100001001000010010000100","0000000010110000101100001011","0000101110101011101010111010","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111000101110001011100010","0000110101001101010011010100","0000111000101110001011100010","0000111111111111111111111111","0000110100001101000011010000","0000101111011011110110111101","0000111000111110001111100011","0000111101101111011011110110","0000111111111111111111111111","0000100111111001111110011111","0000100011001000110010001100","0000011001000110010001100100","0001000000000000000000000000","0000011010100110101001101010","0000100111001001110010011100","0000101000001010000010100000","0000011010110110101101101011","0000011001100110011001100110","0000100000111000001110000011","0000011110110111101101111011","0000100101011001010110010101","0000110001101100011011000110","0000110100001101000011010000","0000110110111101101111011011","0000111000001110000011100000","0000101011001010110010101100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111101101111011011110110","0000111101001111010011110100","0000111110011111100111111001","0000111111111111111111111111","0000011011100110111001101110","0000001101010011010100110101","0000101011001010110010101100","0000110001101100011011000110","0000111011011110110111101101","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111101011111010111110101","0000111111101111111011111110","0000111111011111110111111101","0000101101101011011010110110","0000100100111001001110010011","0000010110010101100101011001","0000001000100010001000100010","0000010100010101000101010001","0000101011101010111010101110","0000100110101001101010011010","0000001000010010000100100001","0000001011010010110100101101","0000110111001101110011011100","0000110010101100101011001010","0000110011111100111111001111","0000110001111100011111000111","0000111110101111101011111010","0000111011101110111011101110","0000111101001111010011110100","0000111111111111111111111111","0000111110011111100111111001","0000100110111001101110011011","0000000100100001001000010010","0000010110100101101001011010","0000011110100111101001111010","0000100011101000111010001110","0000100000111000001110000011","0000100010111000101110001011","0000100101001001010010010100","0000101010011010100110101001","0000110011111100111111001111","0000111010111110101111101011","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111011111110111111101111","0000111011111110111111101111","0000111111011111110111111101","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000100011001000110010001100","0000011111000111110001111100","0000100110011001100110011001","0000010010110100101101001011","0000001010110010101100101011","0000011001100110011001100110","0000010010110100101101001011","0000011110100111101001111010","0000100101011001010110010101","0000011110110111101101111011","0000000101100001011000010110","0000110010001100100011001000","0000111110011111100111111001","0000111111111111111111111111","0000111001001110010011100100","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111010101110101011101010","0000111111111111111111111111","0000111110001111100011111000","0000101100011011000110110001","0000100011101000111010001110","0000001000010010000100100001","0000100000101000001010000010","0000010011000100110001001100","0000101001111010011110100111","0000010000000100000001000000","0000011011110110111101101111","0000011100110111001101110011","0000110101011101010111010101","0000111011101110111011101110","0000111111111111111111111111","0000110101111101011111010111","0000101011111010111110101111","0000100111001001110010011100","0000010000100100001001000010","0000001100100011001000110010","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110111111101111111011111","0000000101000001010000010100","0000010101000101010001010100","0000011010000110100001101000","0000101110011011100110111001","0000101111011011110110111101","0000111000101110001011100010","0000111111001111110011111100","0000111111101111111011111110","0000111110101111101011111010","0000111100001111000011110000","0000111011011110110111101101","0000110011001100110011001100","0000111111011111110111111101","0000110011111100111111001111","0000000110010001100100011001","0000010101000101010001010100","0000111110111111101111111011","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111001101110011011100110","0000111011001110110011101100","0000110100111101001111010011","0000111001101110011011100110","0000111011001110110011101100","0000101100111011001110110011","0000101011011010110110101101","0000111010001110100011101000","0000111101101111011011110110","0000101110111011101110111011","0000100001101000011010000110","0000010101100101011001010110","0000001011010010110100101101","0000011100100111001001110010","0000100000011000000110000001","0000100010001000100010001000","0000011000110110001101100011","0000011111010111110101111101","0000100001001000010010000100","0000011011000110110001101100","0000011100010111000101110001","0000100110101001101010011010","0000110100001101000011010000","0000110111001101110011011100","0000110110101101101011011010","0000111100101111001011110010","0000110110111101101111011011","0000111111111111111111111111","0000111100101111001011110010","0000111101001111010011110100","0000111101111111011111110111","0000111110101111101011111010","0000111110111111101111111011","0000111110101111101011111010","0000111110001111100011111000","0000111101111111011111110111","0000111110011111100111111001","0000110110111101101111011011","0000000010010000100100001001","0000100001001000010010000100","0000100100111001001110010011","0000110010011100100111001001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000111011101110111011101110","0000111100111111001111110011","0000110011111100111111001111","0000101000001010000010100000","0000100000011000000110000001","0001000000000000000000000000","0000011011010110110101101101","0000011110010111100101111001","0000100011111000111110001111","0000010100010101000101010001","0000000000110000001100000011","0000011011010110110101101101","0000101001011010010110100101","0000111000011110000111100001","0000101101111011011110110111","0000111111011111110111111101","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111101101111011011110110","0000111000011110000111100001","0000110011111100111111001111","0000010101110101011101010111","0000001011010010110100101101","0000010111010101110101011101","0000100010011000100110001001","0000101010011010100110101001","0000110100101101001011010010","0000110110101101101011011010","0000111000001110000011100000","0000111001101110011011100110","0000111001001110010011100100","0000110011101100111011001110","0000101110011011100110111001","0000101101111011011110110111","0000100100101001001010010010","0000011100100111001001110010","0000010011010100110101001101","0000010000010100000101000001","0000010101100101011001010110","0000011000000110000001100000","0000001101100011011000110110","0000011011110110111101101111","0000011010000110100001101000","0000000010100000101000001010","0000001001100010011000100110","0000011101110111011101110111","0000101001011010010110100101","0000100001101000011010000110","0000101001111010011110100111","0000010100100101001001010010","0000010100010101000101010001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000111111011111110111111101","0000111110001111100011111000","0000111100001111000011110000","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000110000111100001111000011","0000100000011000000110000001","0000011100100111001001110010","0000001010110010101100101011","0000011110100111101001111010","0000101010111010101110101011","0000010100000101000001010000","0000011111010111110101111101","0000110101111101011111010111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101100001011000010110000","0000100000101000001010000010","0000011101100111011001110110","0000000100110001001100010011","0000110110011101100111011001","0000111111101111111011111110","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000110011011100110111001101","0001000000000000000000000000","0000100101011001010110010101","0000100100001001000010010000","0000110000001100000011000000","0000110111101101111011011110","0000111011101110111011101110","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111101111111011111110111","0000011101110111011101110111","0001000000000000000000000000","0000101100011011000110110001","0000111111101111111011111110","0000111111011111110111111101","0000111110011111100111111001","0000111101011111010111110101","0000111110101111101011111010","0000111010011110100111101001","0000110011001100110011001100","0000110010001100100011001000","0000101010011010100110101001","0000100001011000010110000101","0000110001011100010111000101","0000111111011111110111111101","0000111011111110111111101111","0000100111001001110010011100","0000100001101000011010000110","0001000000000000000000000000","0000011101010111010101110101","0000011111000111110001111100","0000011000110110001101100011","0000010100010101000101010001","0000100110001001100010011000","0000101010101010101010101010","0000111001011110010111100101","0000111011001110110011101100","0000111101101111011011110110","0000111101011111010111110101","0000111110001111100011111000","0000111011001110110011101100","0000111110101111101011111010","0000111100011111000111110001","0000111111001111110011111100","0000111110111111101111111011","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100111111001111110011","0000111011011110110111101101","0000111111111111111111111111","0000011011000110110001101100","0000001001110010011100100111","0000011100010111000101110001","0000100001001000010010000100","0000110111111101111111011111","0000111111001111110011111100","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111000101110001011100010","0000100101011001010110010101","0000011010000110100001101000","0000000010010000100100001001","0000011001110110011101100111","0000100000001000000010000000","0000100010111000101110001011","0000101100101011001010110010","0001000000000000000000000000","0000011001110110011101100111","0000100011011000110110001101","0000101010111010101110101011","0000101011011010110110101101","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111110101111101011111010","0000111100001111000011110000","0000110011011100110111001101","0000100000001000000010000000","0000010001010100010101000101","0000010001010100010101000101","0000001101000011010000110100","0000001001110010011100100111","0000001101100011011000110110","0000001100000011000000110000","0000001000010010000100100001","0000000100100001001000010010","0001000000000000000000000000","0000000011000000110000001100","0000001111100011111000111110","0000001001000010010000100100","0000000101100001011000010110","0000010101000101010001010100","0000010110100101101001011010","0000010110110101101101011011","0000010000110100001101000011","0000001101010011010100110101","0000010110100101101001011010","0000100000111000001110000011","0000001111110011111100111111","0000001011100010111000101110","0000101010111010101110101011","0000100000111000001110000011","0000011010100110101001101010","0000100100111001001110010011","0000000111110001111100011111","0000011110100111101001111010","0000110000101100001011000010","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111011111110111111101","0000111101101111011011110110","0000111110011111100111111001","0000111111001111110011111100","0000110000111100001111000011","0000100111111001111110011111","0000010000100100001001000010","0000000101000001010000010100","0000101100011011000110110001","0000010110110101101101011011","0000011100110111001101110011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111110011111100111111001","0000011111000111110001111100","0000100001001000010010000100","0000000101000001010000010100","0000101100101011001010110010","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000011000000110000001100000","0000000111100001111000011110","0000110111101101111011011110","0000110001101100011011000110","0000101100011011000110110001","0000110001001100010011000100","0000111001111110011111100111","0000111110011111100111111001","0000111110101111101011111010","0000111110001111100011111000","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000100010111000101110001011","0001000000000000000000000000","0000001110110011101100111011","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111110001111100011111000","0000110100001101000011010000","0000101011001010110010101100","0000010101010101010101010101","0000001100110011001100110011","0000100001001000010010000100","0000111001111110011111100111","0000111111111111111111111111","0000100010001000100010001000","0000101100011011000110110001","0000010110100101101001011010","0000001001110010011100100111","0000100001101000011010000110","0000011001010110010101100101","0000011110100111101001111010","0000100111011001110110011101","0000111100011111000111110001","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111010111110101111101011","0000111010001110100011101000","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111100101111001011110010","0000111110101111101011111010","0000111000111110001111100011","0000111110101111101011111010","0000111010101110101011101010","0000101110101011101010111010","0000111100011111000111110001","0000101001111010011110100111","0000000000010000000100000001","0000010001010100010101000101","0000011100110111001101110011","0000100010001000100010001000","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111101011111010111110101","0000011111100111111001111110","0000011010100110101001101010","0001000000000000000000000000","0000010011000100110001001100","0000100100111001001110010011","0000100001001000010010000100","0000100111101001111010011110","0000000111110001111100011111","0000001110100011101000111010","0000101010011010100110101001","0000100000011000000110000001","0000101011001010110010101100","0000111100001111000011110000","0000111101001111010011110100","0000111011011110110111101101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111101111111011111110111","0000110001011100010111000101","0000101010101010101010101010","0000101011001010110010101100","0000100111111001111110011111","0000100000011000000110000001","0000010011100100111001001110","0000001111010011110100111101","0000001010110010101100101011","0000001000010010000100100001","0000000111010001110100011101","0000001010000010100000101000","0000010001110100011101000111","0000011001100110011001100110","0000010110100101101001011010","0000011111100111111001111110","0000011011100110111001101110","0000011000110110001101100011","0000010011000100110001001100","0000001101100011011000110110","0000000101100001011000010110","0000001100000011000000110000","0000000101110001011100010111","0000010001100100011001000110","0000011011010110110101101101","0000101010001010100010101000","0000100000011000000110000001","0000001010010010100100101001","0000001111010011110100111101","0000010110010101100101011001","0000010100100101001001010010","0000101001011010010110100101","0000111110111111101111111011","0000111011011110110111101101","0000111111111111111111111111","0000111010111110101111101011","0000111011011110110111101101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111100111111001111110011","0000111111001111110011111100","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111101111111011111110","0000111001011110010111100101","0000111110011111100111111001","0000110001011100010111000101","0000010000110100001101000011","0000010110010101100101011001","0000011000100110001001100010","0000010111100101111001011110","0000101110111011101110111011","0000111011111110111111101111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000010111000101110001011100","0000001111100011111000111110","0000011010000110100001101000","0000111101001111010011110100","0000111100101111001011110010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000001000010010000100100001","0000010011100100111001001110","0000110110101101101011011010","0000110001101100011011000110","0000111000001110000011100000","0000110001011100010111000101","0000111000011110000111100001","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111010011110100111101001","0000100010111000101110001011","0000000101000001010000010100","0000010010110100101101001011","0000011100010111000101110001","0000111011111110111111101111","0000111101001111010011110100","0000111100101111001011110010","0000111101011111010111110101","0000111111111111111111111111","0000111100101111001011110010","0000110110011101100111011001","0000011110100111101001111010","0000000111000001110000011100","0000000000110000001100000011","0000011111010111110101111101","0000111011101110111011101110","0000111100101111001011110010","0000001011000010110000101100","0000100011001000110010001100","0000000111110001111100011111","0000000111000001110000011100","0000100111101001111010011110","0000010111000101110001011100","0000100001011000010110000101","0000111100011111000111110001","0000110010101100101011001010","0000111110111111101111111011","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111011011110110111101101","0000111011011110110111101101","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000100110111001101110011011","0000110011111100111111001111","0000101110001011100010111000","0000000000100000001000000010","0000001100110011001100110011","0000010011000100110001001100","0000011111100111111001111110","0000110110101101101011011010","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111101111111011111110111","0000011001100110011001100110","0000100010011000100110001001","0000000101100001011000010110","0000001111010011110100111101","0000011111110111111101111111","0000101000011010000110100001","0000011011100110111001101110","0000100000101000001010000010","0001000000000000000000000000","0000101100111011001110110011","0000011100000111000001110000","0000101110001011100010111000","0000110011011100110111001101","0000110010001100100011001000","0000111100011111000111110001","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111100001111000011110000","0000111001101110011011100110","0000110101011101010111010101","0000110010001100100011001000","0000110011101100111011001110","0000110111011101110111011101","0000110011011100110111001101","0000110100111101001111010011","0000110100011101000111010001","0000110010111100101111001011","0000110011111100111111001111","0000110011101100111011001110","0000101100111011001110110011","0000100011111000111110001111","0000011001100110011001100110","0000000110110001101100011011","0000001100010011000100110001","0000000100110001001100010011","0000000010110000101100001011","0000000000100000001000000010","0000001101110011011100110111","0000000000010000000100000001","0000010100010101000101010001","0000010111000101110001011100","0000010111110101111101011111","0000100001001000010010000100","0000100101011001010110010101","0000011100110111001101110011","0000010100100101001001010010","0000001101110011011100110111","0000011011100110111001101110","0000010011000100110001001100","0000101011101010111010101110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100001111000011110000","0000111011101110111011101110","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111001111110011111100111","0000100101001001010010010100","0000001000010010000100100001","0000001001010010010100100101","0000010010010100100101001001","0000011010010110100101101001","0000101010011010100110101001","0000101110111011101110111011","0000110101011101010111010101","0000111111111111111111111111","0000111111101111111011111110","0000110101111101011111010111","0000011100010111000101110001","0000001110000011100000111000","0000000111110001111100011111","0000111111111111111111111111","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111100001111000011110000","0000101010011010100110101001","0001000000000000000000000000","0000101000011010000110100001","0000111101101111011011110110","0000110111111101111111011111","0000111100111111001111110011","0000111001011110010111100101","0000111001001110010011100100","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000110010101100101011001010","0000110011001100110011001100","0000011100010111000101110001","0000011001000110010001100100","0000100101001001010010010100","0000101110011011100110111001","0000111101111111011111110111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000110010011100100111001001","0000010101010101010101010101","0000000010010000100100001001","0000000000110000001100000011","0000110100001101000011010000","0000111111111111111111111111","0000111111001111110011111100","0000100001111000011110000111","0000011100010111000101110001","0000000110110001101100011011","0000001110010011100100111001","0000011110110111101101111011","0000011110110111101101111011","0000101110001011100010111000","0000110100101101001011010010","0000110111011101110111011101","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111100101111001011110010","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000100111101001111010011110","0000101011011010110110101101","0000101110001011100010111000","0000000100010001000100010001","0000001011100010111000101110","0000011100000111000001110000","0000011011110110111101101111","0000101100011011000110110001","0000111110011111100111111001","0000111100111111001111110011","0000111111011111110111111101","0000111101001111010011110100","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000010111000101110001011100","0000101100001011000010110000","0001000000000000000000000000","0000011001000110010001100100","0000100011001000110010001100","0000100100101001001010010010","0000011111100111111001111110","0000011101110111011101110111","0000000000010000000100000001","0000101110011011100110111001","0000011100100111001001110010","0000101001001010010010100100","0000101100111011001110110011","0000110000111100001111000011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000100100011001000110010001","0000011010000110100001101000","0000001100100011001000110010","0000010010100100101001001010","0000001110100011101000111010","0000011111000111110001111100","0000000001110000011100000111","0000000100100001001000010010","0000001100110011001100110011","0000010101100101011001010110","0000011110110111101101111011","0000011101000111010001110100","0000010100110101001101010011","0000011001000110010001100100","0000010100000101000001010000","0000011110100111101001111010","0000010000100100001001000010","0000100011011000110110001101","0000101111111011111110111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111001001110010011100100","0000100011101000111010001110","0000000001100000011000000110","0000001001110010011100100111","0000010011100100111001001110","0000010101000101010001010100","0000100110111001101110011011","0000011110110111101101111011","0000101010011010100110101001","0000111011101110111011101110","0000111011001110110011101100","0000011111000111110001111100","0000010111000101110001011100","0001000000000000000000000000","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111010101110101011101010","0000001111010011110100111101","0000000010100000101000001010","0000110110111101101111011011","0000111111111111111111111111","0000111010101110101011101010","0000110000111100001111000011","0000111111111111111111111111","0000111101101111011011110110","0000111110111111101111111011","0000111010011110100111101001","0000101010001010100010101000","0000011000110110001101100011","0000100011111000111110001111","0000101000111010001110100011","0000111011001110110011101100","0000101111001011110010111100","0000111110101111101011111010","0000111111001111110011111100","0000111111101111111011111110","0000111010101110101011101010","0000111111111111111111111111","0000111110011111100111111001","0000110111011101110111011101","0000100100101001001010010010","0000000101100001011000010110","0000000011010000110100001101","0000001100100011001000110010","0000110001011100010111000101","0000111111011111110111111101","0000111100101111001011110010","0000011110010111100101111001","0000001011110010111100101111","0000010101100101011001010110","0000010001000100010001000100","0000010011110100111101001111","0000100001111000011110000111","0000110010101100101011001010","0000100101011001010110010101","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111111101111111011111110","0000111110011111100111111001","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000100111101001111010011110","0000101100011011000110110001","0000110000111100001111000011","0001000000000000000000000000","0000011000010110000101100001","0000011111100111111001111110","0000100000101000001010000010","0000101101101011011010110110","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000011110100111101001111010","0000010101000101010001010100","0000000100000001000000010000","0000010011110100111101001111","0000100010011000100110001001","0000110000011100000111000001","0000010001010100010101000101","0000011110000111100001111000","0000000001010000010100000101","0000100011011000110110001101","0000100100101001001010010010","0000100010001000100010001000","0000101100001011000010110000","0000110110011101100111011001","0000111110111111101111111011","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111110001111100011111000","0000111011011110110111101101","0000111101001111010011110100","0000111110101111101011111010","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000110011011100110111001101","0000101111111011111110111111","0000101011011010110110101101","0000111100011111000111110001","0000110100111101001111010011","0000101100111011001110110011","0000011111100111111001111110","0000101110111011101110111011","0000101111001011110010111100","0000100000101000001010000010","0001000000000000000000000000","0000000001000000010000000100","0000011011100110111001101110","0000100010101000101010001010","0000101001001010010010100100","0000101010111010101110101011","0000100010001000100010001000","0000100101001001010010010100","0000011111000111110001111100","0000100001111000011110000111","0000100101001001010010010100","0000110010011100100111001001","0000111011001110110011101100","0000111100001111000011110000","0000111100111111001111110011","0000111101111111011111110111","0000111110011111100111111001","0000111110111111101111111011","0000111111011111110111111101","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000100010001000100010001000","0001000000000000000000000000","0000010001000100010001000100","0000010111100101111001011110","0000100000011000000110000001","0000101101011011010110110101","0000100011011000110110001101","0000101111011011110110111101","0000110011101100111011001110","0000100010011000100110001001","0000011011000110110001101100","0000000100010001000100010001","0000101110111011101110111011","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111101111111011111110","0000111111111111111111111111","0000111001111110011111100111","0000110011001100110011001100","0000000010110000101100001011","0000001100000011000000110000","0000111010111110101111101011","0000111010101110101011101010","0000111111011111110111111101","0000110011101100111011001110","0000111111111111111111111111","0000111011111110111111101111","0000110011001100110011001100","0000101110011011100110111001","0000011100100111001001110010","0000100100011001000110010001","0000101001101010011010100110","0000111000001110000011100000","0000111010101110101011101010","0000111010011110100111101001","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101111101011111010111110","0000010111110101111101011111","0001000000000000000000000000","0000001011010010110100101101","0000011001100110011001100110","0000101011011010110110101101","0000111111111111111111111111","0000111100011111000111110001","0000011110110111101101111011","0000010010110100101101001011","0000010100100101001001010010","0001000000000000000000000000","0000010111000101110001011100","0000010111100101111001011110","0000100101101001011010010110","0000110000011100000111000001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111010011110100111101001","0000110000101100001011000010","0000101100101011001010110010","0000101010101010101010101010","0000001001000010010000100100","0000011011110110111101101111","0000011101100111011001110110","0000100001111000011110000111","0000101111111011111110111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000011010010110100101101001","0000001100010011000100110001","0000000001110000011100000111","0000001101110011011100110111","0000101000001010000010100000","0000100100111001001110010011","0000010011000100110001001100","0000100101001001010010010100","0001000000000000000000000000","0000010100000101000001010000","0000011101110111011101110111","0000010011010100110101001101","0000011001010110010101100101","0000100110001001100010011000","0000100111111001111110011111","0000101010001010100010101000","0000101110001011100010111000","0000110010011100100111001001","0000110111011101110111011101","0000111000101110001011100010","0000110101111101011111010111","0000110100011101000111010001","0000111001001110010011100100","0000111111101111111011111110","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111100011111000111110001","0000111111111111111111111111","0000111011001110110011101100","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000110101111101011111010111","0000101001101010011010100110","0000110010101100101011001010","0000111111111111111111111111","0000110101011101010111010101","0000010100100101001001010010","0001000000000000000000000000","0000000100110001001100010011","0000101101101011011010110110","0000110100011101000111010001","0000111111001111110011111100","0000110011101100111011001110","0000111010001110100011101000","0000110000011100000111000001","0000110111111101111111011111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110101011101010111010101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111100001111000011110000","0000111101001111010011110100","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000011101110111011101110111","0000000110000001100000011000","0000010100010101000101010001","0000001101100011011000110110","0000010000000100000001000000","0001000000000000000000000000","0000010101010101010101010101","0000011001010110010101100101","0000010010110100101101001011","0001000000000000000000000000","0001000000000000000000000000","0000011111110111111101111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111100001111000011110000","0000111110101111101011111010","0000111111101111111011111110","0000001101100011011000110110","0000010101110101011101010111","0000011001100110011001100110","0000111101111111011111110111","0000110101001101010011010100","0000111111111111111111111111","0000111111011111110111111101","0000110110101101101011011010","0000110011011100110111001101","0000101011101010111010101110","0000101001001010010010100100","0000110011111100111111001111","0000111100001111000011110000","0000111011001110110011101100","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111100001111000011110000","0000111110001111100011111000","0000101110111011101110111011","0000011110100111101001111010","0000000010000000100000001000","0000000100000001000000010000","0000010011100100111001001110","0000011110010111100101111001","0000101000111010001110100011","0000111011111110111111101111","0000110101101101011011010110","0000101101111011011110110111","0000010010000100100001001000","0000100001111000011110000111","0000010000010100000101000001","0000010111010101110101011101","0000010001110100011101000111","0000011000000110000001100000","0000111011011110110111101101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111000111110001111100011","0000101011011010110110101101","0000101101001011010010110100","0000011000010110000101100001","0000010101010101010101010101","0000100011101000111010001110","0000011000010110000101100001","0000110001111100011111000111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111100011111000111110001","0000111101101111011011110110","0000111110001111100011111000","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000011110100111101001111010","0000000010000000100000001000","0000001010000010100000101000","0000010010010100100101001001","0000100110011001100110011001","0000011101000111010001110100","0000010100110101001101010011","0000011101010111010101110101","0000001001000010010000100100","0000011010010110100101101001","0000011110100111101001111010","0000011111010111110101111101","0000011111100111111001111110","0000100101101001011010010110","0000011101000111010001110100","0000010110110101101101011011","0000100010011000100110001001","0000100010101000101010001010","0000100100101001001010010010","0000101001111010011110100111","0000110001101100011011000110","0000110110011101100111011001","0000110100101101001011010010","0000110000011100000111000001","0000110001011100010111000101","0000110111001101110011011100","0000111101001111010011110100","0000111111001111110011111100","0000111110011111100111111001","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000111011001110110011101100","0000111111111111111111111111","0000111101001111010011110100","0000110010001100100011001000","0000110100101101001011010010","0000111110011111100111111001","0000111111111111111111111111","0000110001111100011111000111","0000010010010100100101001001","0001000000000000000000000000","0000101001101010011010100110","0000100101001001010010010100","0000111010001110100011101000","0000111111111111111111111111","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101011111010111110101","0000111101111111011111110111","0000111111111111111111111111","0000110001101100011011000110","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111100001111000011110000","0000001110010011100100111001","0000001010000010100000101000","0000100001011000010110000101","0000011101010111010101110101","0000101000001010000010100000","0000100111001001110010011100","0000110010101100101011001010","0000011111100111111001111110","0000001100000011000000110000","0000001010010010100100101001","0000000100000001000000010000","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000101101001011010010110100","0000000010010000100100001001","0000101001101010011010100110","0000100101111001011110010111","0000111011101110111011101110","0000110101001101010011010100","0000111100001111000011110000","0000111100111111001111110011","0000110000111100001111000011","0000110011111100111111001111","0000111010011110100111101001","0000111011101110111011101110","0000111111111111111111111111","0000111100111111001111110011","0000111011111110111111101111","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111100001111000011110000","0000111111001111110011111100","0000111111111111111111111111","0000111011011110110111101101","0000110111001101110011011100","0000100010001000100010001000","0000001110110011101100111011","0000000000110000001100000011","0000011111100111111001111110","0000100100111001001110010011","0000011011100110111001101110","0000100101001001010010010100","0000111111111111111111111111","0000111111111111111111111111","0000110100101101001011010010","0001000000000000000000000000","0000011101010111010101110101","0000001010000010100000101000","0000001001110010011100100111","0000010001100100011001000110","0000001101100011011000110110","0000111100011111000111110001","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110011111100111111001111","0000101111111011111110111111","0000100111011001110110011101","0000010010100100101001001010","0000101101111011011110110111","0000010111110101111101011111","0000101111111011111110111111","0000111101001111010011110100","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111101111111011111110111","0000100011101000111010001110","0000000001000000010000000100","0000001101110011011100110111","0000010111110101111101011111","0000011110010111100101111001","0000011000010110000101100001","0000010101000101010001010100","0000001110110011101100111011","0000010111000101110001011100","0000010101010101010101010101","0000001011000010110000101100","0000000111010001110100011101","0000000101000001010000010100","0000000111110001111100011111","0000000011000000110000001100","0001000000000000000000000000","0000000000110000001100000011","0000001001110010011100100111","0000010010010100100101001001","0000010101100101011001010110","0000011000100110001001100010","0000100000011000000110000001","0000101010101010101010101010","0000110001001100010011000100","0000101101001011010010110100","0000101001011010010110100101","0000101011111010111110101111","0000110110111101101111011011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100001111000011110000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000111101011111010111110101","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110001111100011111000","0000111011101110111011101110","0000111100101111001011110010","0000111111111111111111111111","0000111010001110100011101000","0000011110000111100001111000","0000000000110000001100000011","0000011000100110001001100010","0000101001001010010010100100","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111011011110110111101101","0000111000101110001011100010","0000110111101101111011011110","0000111001011110010111100101","0000111010111110101111101011","0000111011111110111111101111","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000110100111101001111010011","0000101111101011111010111110","0000111000001110000011100000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000101110011011100110111001","0000000011100000111000001110","0000010100110101001101010011","0000100011111000111110001111","0000101111001011110010111100","0000110011101100111011001110","0000111111111111111111111111","0000110000101100001011000010","0000100110111001101110011011","0000011100100111001001110010","0001000000000000000000000000","0000111011101110111011101110","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000000101010001010100010101","0000100101001001010010010100","0000101001011010010110100101","0000101010111010101110101011","0000110010111100101111001011","0000111010101110101011101010","0000111111001111110011111100","0000111101101111011011110110","0000111110001111100011111000","0000111100011111000111110001","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111111111111111111111111","0000111100011111000111110001","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111101111111011111110111","0000111110011111100111111001","0000111110101111101011111010","0000111010001110100011101000","0000101001001010010010100100","0000100101111001011110010111","0001000000000000000000000000","0000001110010011100100111001","0000110000001100000011000000","0000101101101011011010110110","0000011100010111000101110001","0000101100101011001010110010","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000011010010110100101101001","0000011010010110100101101001","0000010111010101110101011101","0001000000000000000000000000","0000001100110011001100110011","0000000001100000011000000110","0000111111111111111111111111","0000111011001110110011101100","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000110110001101100011011000","0000101010001010100010101000","0000100100101001001010010010","0000001101110011011100110111","0000010111000101110001011100","0000100101011001010110010101","0000101110001011100010111000","0000111100011111000111110001","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111011011110110111101101","0000111101011111010111110101","0000111110111111101111111011","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111101011111010111110101","0000011101100111011001110110","0000001110010011100100111001","0000000110110001101100011011","0000010010010100100101001001","0000011000100110001001100010","0000010001000100010001000100","0000010101010101010101010101","0000010001010100010101000101","0000000010010000100100001001","0000000001100000011000000110","0000010000010100000101000001","0000010100100101001001010010","0000100000011000000110000001","0000100101001001010010010100","0000100110011001100110011001","0000101001111010011110100111","0000101011001010110010101100","0000011100110111001101110011","0000010001000100010001000100","0000001110000011100000111000","0000001100000011000000110000","0000001010010010100100101001","0000010001010100010101000101","0000011100100111001001110010","0000100001111000011110000111","0000100001011000010110000101","0000100001111000011110000111","0000101000001010000010100000","0000110100001101000011010000","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000101100011011000110110001","0000100001111000011110000111","0000000001100000011000000110","0000010010000100100001001000","0000101000011010000110100001","0000111101111111011111110111","0000111101001111010011110100","0000111011111110111111101111","0000110001101100011011000110","0000101010011010100110101001","0000100010001000100010001000","0000011010010110100101101001","0000011000100110001001100010","0000011100100111001001110010","0000100110001001100010011000","0000110011111100111111001111","0000111111011111110111111101","0000111100101111001011110010","0000111010001110100011101000","0000100011101000111010001110","0000110011001100110011001100","0000111011111110111111101111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000110111111101111111011111","0000110111011101110111011101","0000000101110001011100010111","0000000111000001110000011100","0000100010001000100010001000","0000110010111100101111001011","0000111111101111111011111110","0000111111001111110011111100","0000111000111110001111100011","0000100010101000101010001010","0000010111100101111001011110","0000010000110100001101000011","0000111000001110000011100000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000101000001010000010100000","0000000100010001000100010001","0000111111111111111111111111","0000100000101000001010000010","0000110001001100010011000100","0000101000011010000110100001","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111101001111010011110100","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111100001111000011110000","0000111101101111011011110110","0000111111011111110111111101","0000111110001111100011111000","0000111101001111010011110100","0000111101101111011011110110","0000111111101111111011111110","0000110100101101001011010010","0000110010111100101111001011","0000110111011101110111011101","0000010101100101011001010110","0000000001110000011100000111","0000001110110011101100111011","0000111001011110010111100101","0000101011101010111010101110","0000011000110110001101100011","0000110101011101010111010101","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000101111011011110110111101","0000011110010111100101111001","0000001110100011101000111010","0000000100010001000100010001","0000001111000011110000111100","0000000000100000001000000010","0000111011011110110111101101","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111111101111111011111110","0000111110111111101111111011","0000101110111011101110111011","0000011011010110110101101101","0000010000110100001101000011","0000001110000011100000111000","0000011000110110001101100011","0000101000011010000110100001","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000111100011111000111110001","0000111100011111000111110001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111110001111100011111000","0000111110001111100011111000","0000111101011111010111110101","0000101100101011001010110010","0000010100110101001101010011","0000001011110010111100101111","0000000100010001000100010001","0000010101000101010001010100","0000010100010101000101010001","0000010001000100010001000100","0000010100010101000101010001","0000000000110000001100000011","0000011100110111001101110011","0000100000011000000110000001","0000011110010111100101111001","0000011000000110000001100000","0000100000011000000110000001","0000100111101001111010011110","0000100110001001100010011000","0000101110101011101010111010","0000110000111100001111000011","0000111000111110001111100011","0000110100001101000011010000","0000101100011011000110110001","0000110100001101000011010000","0000111001011110010111100101","0000101001001010010010100100","0000010011110100111101001111","0000000111010001110100011101","0000001100100011001000110010","0000010000010100000101000001","0000100010101000101010001010","0000101000101010001010100010","0000110010011100100111001001","0000111011111110111111101111","0000111111111111111111111111","0000111101011111010111110101","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111011111110111111101111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000101101101011011010110110","0000010111010101110101011101","0001000000000000000000000000","0000011001100110011001100110","0000100000011000000110000001","0000101101111011011110110111","0000101001001010010010100100","0000100000001000000010000000","0000011111110111111101111111","0000010110100101101001011010","0000001101110011011100110111","0000000010000000100000001000","0000000000010000000100000001","0000001100110011001100110011","0000011110010111100101111001","0000110001001100010011000100","0000111101101111011011110110","0000101010001010100010101000","0000101001111010011110100111","0000101101111011011110110111","0000111100101111001011110010","0000110101111101011111010111","0000111101111111011111110111","0000111111101111111011111110","0000111101101111011011110110","0000111101011111010111110101","0000110110011101100111011001","0000110111111101111111011111","0000011000100110001001100010","0001000000000000000000000000","0000011100110111001101110011","0000110111001101110011011100","0000111111101111111011111110","0000111111001111110011111100","0000110011001100110011001100","0000100100011001000110010001","0000010111010101110101011101","0000001111110011111100111111","0000101101111011011110110111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111110001111100011111000","0000110101111101011111010111","0000111111111111111111111111","0000110111111101111111011111","0001000000000000000000000000","0000111011011110110111101101","0000111010001110100011101000","0000011111110111111101111111","0000111000111110001111100011","0000100110011001100110011001","0000111111111111111111111111","0000111100001111000011110000","0000111010101110101011101010","0000111010111110101111101011","0000111111111111111111111111","0000111011101110111011101110","0000111110111111101111111011","0000111111111111111111111111","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000101111111011111110111111","0000111010101110101011101010","0000100111001001110010011100","0000100001101000011010000110","0000001101110011011100110111","0000001011100010111000101110","0000100000101000001010000010","0000111001011110010111100101","0000101111001011110010111100","0000100011111000111110001111","0000111110101111101011111010","0000111101011111010111110101","0000111110111111101111111011","0000111101111111011111110111","0000111011111110111111101111","0000011110010111100101111001","0000101001111010011110100111","0000000011010000110100001101","0000000111110001111100011111","0001000000000000000000000000","0000101011111010111110101111","0000111001001110010011100100","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111011111110111111101111","0000101100001011000010110000","0000001011100010111000101110","0000100001101000011010000110","0000011011000110110001101100","0000011101110111011101110111","0000111110011111100111111001","0000111101111111011111110111","0000111100111111001111110011","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111110101111101011111010","0000111110111111101111111011","0000111111101111111011111110","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000101111101011111010111110","0000100110011001100110011001","0000000101100001011000010110","0000001110100011101000111010","0000001001100010011000100110","0000001110110011101100111011","0000010101100101011001010110","0000010101010101010101010101","0000000101100001011000010110","0000100100011001000110010001","0000100001101000011010000110","0000101101011011010110110101","0000110000101100001011000010","0000110101001101010011010100","0000111111001111110011111100","0000111111111111111111111111","0000111100101111001011110010","0000111101101111011011110110","0000111111101111111011111110","0000111011111110111111101111","0000111101001111010011110100","0000111010101110101011101010","0000110100001101000011010000","0000111000111110001111100011","0000111111001111110011111100","0000111011001110110011101100","0000111011111110111111101111","0000110001111100011111000111","0000100010111000101110001011","0000100101011001010110010101","0000100111001001110010011100","0000101110011011100110111001","0000110101101101011011010110","0000111110111111101111111011","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111101111111011111110111","0000111110011111100111111001","0000111111011111110111111101","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111100101111001011110010","0000111110011111100111111001","0000101111001011110010111100","0000001101100011011000110110","0000000011000000110000001100","0000011110000111100001111000","0000011001000110010001100100","0000100101001001010010010100","0000100100001001000010010000","0000001000000010000000100000","0000000111000001110000011100","0000100110011001100110011001","0000110000001100000011000000","0000101111011011110110111101","0000100011111000111110001111","0000000001010000010100000101","0001000000000000000000000000","0000101100111011001110110011","0000101110111011101110111011","0000110000111100001111000011","0000101000011010000110100001","0000111111111111111111111111","0000101011111010111110101111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000110100111101001111010011","0000110011001100110011001100","0000011110000111100001111000","0000000100100001001000010010","0000000111000001110000011100","0000110010001100100011001000","0000111111101111111011111110","0000111110111111101111111011","0000111001011110010111100101","0000100111001001110010011100","0000011010010110100101101001","0000011100100111001001110010","0000100111101001111010011110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111100011111000111110001","0000111101011111010111110101","0000111111111111111111111111","0000111011011110110111101101","0000010001110100011101000111","0000100111101001111010011110","0000111101101111011011110110","0000110000001100000011000000","0000100111001001110010011100","0000101100011011000110110001","0000101111111011111110111111","0000111000001110000011100000","0000111111111111111111111111","0000111101011111010111110101","0000110101111101011111010111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111101111111011111110111","0000110001111100011111000111","0000110010011100100111001001","0000100001001000010010000100","0000101101101011011010110110","0000100011101000111010001110","0000000011100000111000001110","0000011100100111001001110010","0000011101110111011101110111","0000111011011110110111101101","0000110110001101100011011000","0000100111101001111010011110","0000111111111111111111111111","0000111100011111000111110001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000100101001001010010010100","0000110100011101000111010001","0000100110001001100010011000","0000000000110000001100000011","0000010001110100011101000111","0000001111010011110100111101","0000110000101100001011000010","0000111111111111111111111111","0000111100101111001011110010","0000111101011111010111110101","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000110111001101110011011100","0000010010100100101001001010","0000011000110110001101100011","0000010001010100010101000101","0000100011001000110010001100","0000110100101101001011010010","0000111110001111100011111000","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111101101111011011110110","0000111110101111101011111010","0000111111101111111011111110","0000111111011111110111111101","0000111110101111101011111010","0000111111101111111011111110","0000111110011111100111111001","0000111111011111110111111101","0000111110011111100111111001","0000111110111111101111111011","0000111000001110000011100000","0000100110101001101010011010","0000011010010110100101101001","0001000000000000000000000000","0000010101010101010101010101","0001000000000000000000000000","0000010000010100000101000001","0000001101000011010000110100","0000001010000010100000101000","0000100110101001101010011010","0000100111011001110110011101","0000110101101101011011010110","0000111110001111100011111000","0000111000111110001111100011","0000111010101110101011101010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111000101110001011100010","0000101111111011111110111111","0000101001111010011110100111","0000101101011011010110110101","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111010111110101111101011","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000011111000111110001111100","0000001100110011001100110011","0000010000110100001101000011","0000100101001001010010010100","0000100101101001011010010110","0000000100000001000000010000","0000100010011000100110001001","0000111011001110110011101100","0000111001101110011011100110","0000111100001111000011110000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000100100001001000010010000","0001000000000000000000000000","0000001101010011010100110101","0000100001011000010110000101","0000001001100010011000100110","0000110000111100001111000011","0000110111001101110011011100","0000110110111101101111011011","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000110101111101011111010111","0000100111001001110010011100","0000011100010111000101110001","0000001101110011011100110111","0000000000010000000100000001","0000100100111001001110010011","0000111011101110111011101110","0000111111111111111111111111","0000111111101111111011111110","0000101000101010001010100010","0000100100111001001110010011","0000010111110101111101011111","0000011010100110101001101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111110011111100111111001","0000111111011111110111111101","0000111100101111001011110010","0000101010111010101110101011","0000001010110010101100101011","0000111110101111101011111010","0000111110101111101011111010","0000101000111010001110100011","0000101001111010011110100111","0000101100111011001110110011","0000110001001100010011000100","0000101101001011010010110100","0000111100001111000011110000","0000111111111111111111111111","0000101011101010111010101110","0000111010111110101111101011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000101101111011011110110111","0000110110111101101111011011","0000101001101010011010100110","0000111011101110111011101110","0000100110111001101110011011","0000000001010000010100000101","0000100110101001101010011010","0000100100011001000110010001","0000011010010110100101101001","0000111100101111001011110010","0000111000111110001111100011","0000101100111011001110110011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000110110101101101011011010","0000101111111011111110111111","0000111010001110100011101000","0001000000000000000000000000","0000000000100000001000000010","0000010100110101001101010011","0000100000101000001010000010","0000111001011110010111100101","0000111111111111111111111111","0000111100001111000011110000","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111110011111100111111001","0000110100001101000011010000","0000010011110100111101001111","0000101011101010111010101110","0000010001010100010101000101","0000101010001010100010101000","0000111111111111111111111111","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111100111111001111110011","0000100100111001001110010011","0000011101010111010101110101","0000010000110100001101000011","0000000100110001001100010011","0000010111110101111101011111","0001000000000000000000000000","0000001001010010010100100101","0000000001010000010100000101","0000100100001001000010010000","0000100000011000000110000001","0000110011101100111011001110","0000111101111111011111110111","0000111111111111111111111111","0000111100011111000111110001","0000111011101110111011101110","0000111110011111100111111001","0000111101001111010011110100","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111101001111010011110100","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111010011110100111101001","0000101110101011101010111010","0000101001011010010110100101","0000111100101111001011110010","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111100001111000011110000","0000111100001111000011110000","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111101011111010111110101","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111011101110111011101110","0000111111001111110011111100","0000111100011111000111110001","0000011100110111001101110011","0001000000000000000000000000","0000110001011100010111000101","0000000000100000001000000010","0000011010000110100001101000","0000110010011100100111001001","0000110011001100110011001100","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000101111011011110110111101","0001000000000000000000000000","0000001111010011110100111101","0000100100011001000110010001","0000100001011000010110000101","0000101001111010011110100111","0000110110011101100111011001","0000111101011111010111110101","0000111111101111111011111110","0000111101101111011011110110","0000111010011110100111101001","0000100001011000010110000101","0000011010010110100101101001","0000011000110110001101100011","0000001001000010010000100100","0000000001010000010100000101","0000111011011110110111101101","0000111001111110011111100111","0000111111111111111111111111","0000110110111101101111011011","0000100100101001001010010010","0000001111000011110000111100","0000000111000001110000011100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110101101101011011010","0000000110110001101100011011","0000101110101011101010111010","0000111111101111111011111110","0000111111011111110111111101","0000011001010110010101100101","0000101011011010110110101101","0000110001001100010011000100","0000111001001110010011100100","0000101011001010110010101100","0000111111111111111111111111","0000111100111111001111110011","0000111011001110110011101100","0000110000111100001111000011","0000110111111101111111011111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111101001111010011110100","0000101110001011100010111000","0000101110111011101110111011","0000110001001100010011000100","0000111000001110000011100000","0000111010111110101111101011","0000100000101000001010000010","0000000000100000001000000010","0000011000000110000001100000","0000100101011001010110010101","0000101101011011010110110101","0000101000111010001110100011","0000111111011111110111111101","0000110111111101111111011111","0000111010001110100011101000","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111101001111010011110100","0000111111111111111111111111","0000110111011101110111011101","0000101011001010110010101100","0000011101010111010101110101","0001000000000000000000000000","0000001000100010001000100010","0000010110100101101001011010","0000111011011110110111101101","0000111110001111100011111000","0000111110111111101111111011","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111110011111100111111001","0000110100001101000011010000","0000100001001000010010000100","0000100101001001010010010100","0000011011000110110001101100","0000110101011101010111010101","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000101010001010100010101000","0000100100011001000110010001","0000011001000110010001100100","0000000010010000100100001001","0000010101110101011101010111","0000011010010110100101101001","0000000100010001000100010001","0000000101010001010100010101","0000010100000101000001010000","0000011101110111011101110111","0000100110111001101110011011","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000110101011101010111010101","0000101101001011010010110100","0000111010101110101011101010","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111111001111110011111100","0000111111101111111011111110","0000111101011111010111110101","0000110111111101111111011111","0000110011011100110111001101","0000111010101110101011101010","0000110000111100001111000011","0000111101001111010011110100","0000110111001101110011011100","0000111010111110101111101011","0000110101101101011011010110","0000111100011111000111110001","0000111111111111111111111111","0000110100111101001111010011","0000111111111111111111111111","0000111100001111000011110000","0000101010001010100010101000","0000000010110000101100001011","0000001011100010111000101110","0000010011110100111101001111","0000101110101011101010111010","0000110000001100000011000000","0000111111011111110111111101","0000111110001111100011111000","0000111110001111100011111000","0000111011011110110111101101","0000111010011110100111101001","0000111111111111111111111111","0000111010001110100011101000","0000110010101100101011001010","0000101001011010010110100101","0000000000010000000100000001","0000001011010010110100101101","0000011010000110100001101000","0000011100100111001001110010","0000110111111101111111011111","0000111011111110111111101111","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000101000001010000010100000","0000010011110100111101001111","0000010011110100111101001111","0000010111010101110101011101","0000000011010000110100001101","0000011001100110011001100110","0000111111111111111111111111","0000111110101111101011111010","0000111010001110100011101000","0000100101101001011010010110","0000001101010011010100110101","0000000000110000001100000011","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000100101001001010010010100","0000011000100110001001100010","0000111111111111111111111111","0000111111111111111111111111","0000101111111011111110111111","0000010101000101010001010100","0000100000011000000110000001","0000101011101010111010101110","0000111011001110110011101100","0000101011111010111110101111","0000111010101110101011101010","0000111111111111111111111111","0000111110011111100111111001","0000111000011110000111100001","0000110100101101001011010010","0000111001101110011011100110","0000111100101111001011110010","0000110010101100101011001010","0000011101100111011001110110","0000100001011000010110000101","0000100100111001001110010011","0000101111011011110110111101","0000111111111111111111111111","0000101111111011111110111111","0000100000111000001110000011","0000001011000010110000101100","0000100111111001111110011111","0000110010101100101011001010","0000101110001011100010111000","0000110101011101010111010101","0000111111111111111111111111","0000111010101110101011101010","0000111111101111111011111110","0000111100101111001011110010","0000111111101111111011111110","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000100100001001000010010000","0000000100010001000100010001","0000001011100010111000101110","0000001110010011100100111001","0000100111011001110110011101","0000111011101110111011101110","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000110111001101110011011100","0000100011111000111110001111","0000100011011000110110001101","0000011111100111111001111110","0000111101101111011011110110","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111100101111001011110010","0000111011001110110011101100","0000111011011110110111101101","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110110101101101011011010","0000100110101001101010011010","0000010100010101000101010001","0000101100111011001110110011","0000010010010100100101001001","0000000000110000001100000011","0000100001101000011010000110","0000010110010101100101011001","0001000000000000000000000000","0000001110110011101100111011","0000010101110101011101010111","0000010101110101011101010111","0000110110111101101111011011","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000111100101111001011110010","0000111100101111001011110010","0000111110101111101011111010","0000111011101110111011101110","0000111111111111111111111111","0000111011111110111111101111","0000111100011111000111110001","0000111110011111100111111001","0000111111011111110111111101","0000111110001111100011111000","0000111110001111100011111000","0000111110011111100111111001","0000111101011111010111110101","0000111101001111010011110100","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100011101000111010001","0000110011001100110011001100","0000111111001111110011111100","0000111111011111110111111101","0000111110001111100011111000","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111000101110001011100010","0000110110001101100011011000","0000111001011110010111100101","0000101110001011100010111000","0000111111111111111111111111","0000101101001011010010110100","0000110001001100010011000100","0000111111011111110111111101","0000111111001111110011111100","0000101110101011101010111010","0000111101001111010011110100","0000111110011111100111111001","0000101101111011011110110111","0000001010100010101000101010","0001000000000000000000000000","0000101111011011110110111101","0000100101111001011110010111","0000111100101111001011110010","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000110011111100111111001111","0000110000001100000011000000","0000010010100100101001001010","0001000000000000000000000000","0000010111010101110101011101","0000010111100101111001011110","0000100110011001100110011001","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111000001110000011100000","0000011100010111000101110001","0000010000010100000101000001","0000011101110111011101110111","0000011010010110100101101001","0000000001010000010100000101","0000101101101011011010110110","0000111111111111111111111111","0000111000011110000111100001","0000101010001010100010101000","0000000110000001100000011000","0000000011100000111000001110","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110110111101101111011011","0000010000000100000001000000","0000111000111110001111100011","0000111111011111110111111101","0000111010011110100111101001","0000100000001000000010000000","0000010111010101110101011101","0000100101101001011010010110","0000100000011000000110000001","0000101110011011100110111001","0000100110011001100110011001","0000111100001111000011110000","0000111110001111100011111000","0000111111111111111111111111","0000111010011110100111101001","0000110111001101110011011100","0000101010101010101010101010","0000011111110111111101111111","0000100000011000000110000001","0000100001011000010110000101","0000100011111000111110001111","0000100010011000100110001001","0000101100111011001110110011","0000101001111010011110100111","0000110001001100010011000100","0000010101100101011001010110","0000110000011100000111000001","0000100011011000110110001101","0000111101101111011011110110","0000111010101110101011101010","0000101110011011100110111001","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000111100101111001011110010","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000110111111101111111011111","0000111010001110100011101000","0000111110101111101011111010","0000111001001110010011100100","0000000001100000011000000110","0000000111110001111100011111","0000001001100010011000100110","0000010111000101110001011100","0000111011111110111111101111","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111011111110111111101111","0000101111101011111010111110","0000110000101100001011000010","0000110010111100101111001011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000110010111100101111001011","0000110001001100010011000100","0000111000101110001011100010","0000111111111111111111111111","0000111101011111010111110101","0000100100111001001110010011","0000011001000110010001100100","0000011000100110001001100010","0000010011010100110101001101","0000011011110110111101101111","0000000010010000100100001001","0000010110000101100001011000","0000100000011000000110000001","0000011000010110000101100001","0000000000010000000100000001","0000000011000000110000001100","0000011101110111011101110111","0000010001010100010101000101","0000111001101110011011100110","0000111000011110000111100001","0000111110111111101111111011","0000111100101111001011110010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000111100011111000111110001","0000110010111100101111001011","0000111000011110000111100001","0000111110001111100011111000","0000111101011111010111110101","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000110010101100101011001010","0000110111111101111111011111","0000110000111100001111000011","0000101000101010001010100010","0000100100101001001010010010","0000111111111111111111111111","0000110100001101000011010000","0000101110101011101010111010","0000111111111111111111111111","0000111111001111110011111100","0000110000011100000111000001","0000001100110011001100110011","0000000000100000001000000010","0000100001001000010010000100","0000101111011011110110111101","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111110111111101111111011","0000111110001111100011111000","0000111101001111010011110100","0000111010111110101111101011","0000111100111111001111110011","0000111111111111111111111111","0000101001001010010010100100","0000101000011010000110100001","0000001100010011000100110001","0000010001100100011001000110","0000011111010111110101111101","0000100000111000001110000011","0000110111111101111111011111","0000111101111111011111110111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000110000111100001111000011","0000011010000110100001101000","0000011110110111101101111011","0000011001000110010001100100","0000011000000110000001100000","0001000000000000000000000000","0000110011001100110011001100","0000111001001110010011100100","0000100010111000101110001011","0000000100010001000100010001","0000000110110001101100011011","0000100110001001100010011000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000110000001100000011000000","0000010111010101110101011101","0000111010101110101011101010","0000110100011101000111010001","0000111101011111010111110101","0000100011111000111110001111","0000001110110011101100111011","0000011101010111010101110101","0000100010111000101110001011","0000010001000100010001000100","0000100001101000011010000110","0000101011001010110010101100","0000100110101001101010011010","0000100110111001101110011011","0000100011011000110110001101","0000001110110011101100111011","0000000011000000110000001100","0000000010000000100000001000","0001000000000000000000000000","0000000010110000101100001011","0000001011010010110100101101","0000010000100100001001000010","0000101101011011010110110101","0000101000011010000110100001","0000100101011001010110010101","0000110100101101001011010010","0000100111011001110110011101","0000111001001110010011100100","0000110111011101110111011101","0000110001001100010011000100","0000101111101011111010111110","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100111111001111110011","0000111101101111011011110110","0000110001001100010011000100","0000111011111110111111101111","0000111101001111010011110100","0000011110010111100101111001","0000000101000001010000010100","0000011000100110001001100010","0000010001010100010101000101","0000110101011101010111010101","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111111101111111011111110","0000111110111111101111111011","0000110000101100001011000010","0000110111011101110111011101","0000110110011101100111011001","0000111100111111001111110011","0000111101101111011011110110","0000111111111111111111111111","0000111111001111110011111100","0000111100101111001011110010","0000111110111111101111111011","0000111101101111011011110110","0000111100011111000111110001","0000111100001111000011110000","0000111011101110111011101110","0000111000001110000011100000","0000110010101100101011001010","0000101110001011100010111000","0000011110100111101001111010","0000010011010100110101001101","0000010001110100011101000111","0000010010000100100001001000","0000010100110101001101010011","0000000111100001111000011110","0001000000000000000000000000","0000100001101000011010000110","0000100001001000010010000100","0000011000000110000001100000","0000000110100001101000011010","0000000101100001011000010110","0000010111110101111101011111","0000011000110110001101100011","0000101110111011101110111011","0000111100011111000111110001","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111110101111101011111010","0000111111111111111111111111","0000111011111110111111101111","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000110100101101001011010010","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111000101110001011100010","0000110111001101110011011100","0000111001101110011011100110","0000111100111111001111110011","0000110010111100101111001011","0000110110111101101111011011","0000101101101011011010110110","0000101111111011111110111111","0000010111000101110001011100","0000011101100111011001110110","0000111010101110101011101010","0000100110111001101110011011","0000110110011101100111011001","0000111111111111111111111111","0000111100011111000111110001","0000111000111110001111100011","0000000010010000100100001001","0001000000000000000000000000","0000011111010111110101111101","0000101110011011100110111001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000011010100110101001101010","0000010111110101111101011111","0000001100010011000100110001","0000011100000111000001110000","0000101110001011100010111000","0000101101011011010110110101","0000110111101101111011011110","0000111110111111101111111011","0000111111111111111111111111","0000111011011110110111101101","0000101110001011100010111000","0000011000110110001101100011","0000101010001010100010101000","0000100101001001010010010100","0000011110000111100001111000","0000010101010101010101010101","0000001011010010110100101101","0000100101001001010010010100","0000011110110111101101111011","0000001110010011100100111001","0000010100000101000001010000","0000000001010000010100000101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101111111011111110111","0000001011110010111100101111","0000101000101010001010100010","0000110001011100010111000101","0000101101001011010010110100","0000110100011101000111010001","0000101100111011001110110011","0000100101101001011010010110","0000001110110011101100111011","0000011001110110011101100111","0000001101110011011100110111","0000000011010000110100001101","0000010101000101010001010100","0000011001110110011101100111","0000010010110100101101001011","0000000101000001010000010100","0000001010010010100100101001","0000010001110100011101000111","0000001101110011011100110111","0000010001110100011101000111","0000010111110101111101011111","0000010010110100101101001011","0000011011000110110001101100","0000000001000000010000000100","0000000001010000010100000101","0000100110001001100010011000","0000101111101011111010111110","0000011101110111011101110111","0000101001001010010010100100","0000110010101100101011001010","0000110110001101100011011000","0000110110101101101011011010","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000101010111010101110101011","0000111101111111011111110111","0000011010000110100001101000","0001000000000000000000000000","0000010010010100100101001001","0000010001010100010101000101","0000101000111010001110100011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000101010111010101110101011","0000111111111111111111111111","0000101000001010000010100000","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000111111011111110111111101","0000111101111111011111110111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000101110101011101010111010","0000110100011101000111010001","0000101111011011110110111101","0000010110000101100001011000","0000010010110100101101001011","0000010001110100011101000111","0000000111010001110100011101","0001000000000000000000000000","0000001110100011101000111010","0000100000111000001110000011","0000100000011000000110000001","0000011101000111010001110100","0000100011001000110010001100","0000000001110000011100000111","0001000000000000000000000000","0000010110010101100101011001","0000010010100100101001001010","0000100111011001110110011101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111101111111011111110111","0000111100011111000111110001","0000111111101111111011111110","0000111110101111101011111010","0000111100001111000011110000","0000111111101111111011111110","0000111110101111101011111010","0000111110101111101011111010","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111110111111101111111011","0000111011011110110111101101","0000111101111111011111110111","0000111101001111010011110100","0000111100011111000111110001","0000111100001111000011110000","0000110001011100010111000101","0000111111111111111111111111","0000111100111111001111110011","0000111101111111011111110111","0000110110111101101111011011","0000111010001110100011101000","0000101110011011100110111001","0000101111101011111010111110","0000011011100110111001101110","0000011111100111111001111110","0000010101000101010001010100","0000100010011000100110001001","0000101010001010100010101000","0000100010011000100110001001","0000111000011110000111100001","0000111111111111111111111111","0000111110101111101011111010","0000111001101110011011100110","0000000001100000011000000110","0000010001110100011101000111","0000010010100100101001001010","0000110101011101010111010101","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000010111110101111101011111","0000010010100100101001001010","0000010111010101110101011101","0000010110010101100101011001","0000110110111101101111011011","0000111011111110111111101111","0000101010001010100010101000","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000110011001100110011001100","0000100000001000000010000000","0000100000001000000010000000","0000101100011011000110110001","0000110100011101000111010001","0000001111110011111100111111","0000010001000100010001000100","0000010111110101111101011111","0000001010110010101100101011","0000001111000011110000111100","0000010110000101100001011000","0000000000100000001000000010","0000100010101000101010001010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111101001111010011110100","0000111110101111101011111010","0000111111111111111111111111","0000111010101110101011101010","0000110100111101001111010011","0000000000010000000100000001","0000110001111100011111000111","0000100101001001010010010100","0000100110101001101010011010","0000100101111001011110010111","0000110110111101101111011011","0000110100011101000111010001","0000011110100111101001111010","0000011101010111010101110101","0000010000000100000001000000","0000001110010011100100111001","0000010100010101000101010001","0000110010011100100111001001","0000101101101011011010110110","0000011011000110110001101100","0000011010010110100101101001","0000000010000000100000001000","0000000100110001001100010011","0000000100010001000100010001","0000001010000010100000101000","0001000000000000000000000000","0000000101010001010100010101","0000000111110001111100011111","0000100000011000000110000001","0000101101101011011010110110","0000101010011010100110101001","0000110011011100110111001101","0000111001111110011111100111","0000111011111110111111101111","0000111001011110010111100101","0000111011101110111011101110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111110111111101111111011","0000111110111111101111111011","0000111010101110101011101010","0000110100111101001111010011","0000101011111010111110101111","0000000110000001100000011000","0000000001100000011000000110","0000001000100010001000100010","0000001111100011111000111110","0000100000111000001110000011","0000111101001111010011110100","0000111111011111110111111101","0000111110001111100011111000","0000111101101111011011110110","0000111100111111001111110011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000110000111100001111000011","0000111111111111111111111111","0000111000001110000011100000","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111101111111011111110111","0000111110011111100111111001","0000111100011111000111110001","0000101100011011000110110001","0000100000101000001010000010","0000001101010011010100110101","0000000000100000001000000010","0000001101100011011000110110","0000100000011000000110000001","0000011111100111111001111110","0000100011101000111010001110","0000011111110111111101111111","0000010111000101110001011100","0000100001111000011110000111","0001000000000000000000000000","0000010001010100010101000101","0000010000100100001001000010","0000011000110110001101100011","0000101010001010100010101000","0000110110111101101111011011","0000110101101101011011010110","0000111010011110100111101001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111011111110111111101111","0000110110101101101011011010","0000111001001110010011100100","0000110100001101000011010000","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111000001110000011100000","0000110110101101101011011010","0000111111111111111111111111","0000110111111101111111011111","0000111111111111111111111111","0000111011101110111011101110","0000101100111011001110110011","0000110110001101100011011000","0000111001111110011111100111","0000110000101100001011000010","0000100111111001111110011111","0000100110101001101010011010","0000100011101000111010001110","0000100000101000001010000010","0000011001010110010101100101","0000001111100011111000111110","0000010110010101100101011001","0000011110110111101101111011","0000110011011100110111001101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000101001111010011110100111","0000100000011000000110000001","0000000100100001001000010010","0000001010100010101000101010","0000110111001101110011011100","0000111110111111101111111011","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000011000010110000101100001","0000001100100011001000110010","0000101001101010011010100110","0000100011011000110110001101","0000110110001101100011011000","0000111111101111111011111110","0000111111001111110011111100","0000110111011101110111011101","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000101101001011010010110100","0000011110110111101101111011","0000100000001000000010000000","0000111100111111001111110011","0000110010111100101111001011","0000100110001001100010011000","0000100110011001100110011001","0000010101010101010101010101","0000000000010000000100000001","0000010101110101011101010111","0000001101010011010100110101","0000001100110011001100110011","0000111101101111011011110110","0000111011001110110011101100","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000011110010111100101111001","0000001010010010100100101001","0000110101001101010011010100","0000100111111001111110011111","0000101110111011101110111011","0000101110001011100010111000","0000110110101101101011011010","0000111000001110000011100000","0000100100111001001110010011","0000110000001100000011000000","0000010000110100001101000011","0000001011010010110100101101","0000000111000001110000011100","0000011001010110010101100101","0000010101110101011101010111","0000100001011000010110000101","0000011011000110110001101100","0000101100001011000010110000","0000110000011100000111000001","0000100010011000100110001001","0000101101111011011110110111","0000110111001101110011011100","0000101010111010101110101011","0000001010000010100000101000","0000100000011000000110000001","0000101110001011100010111000","0000011111000111110001111100","0000111100001111000011110000","0000111111001111110011111100","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111110001111100011111000","0000111110001111100011111000","0000111101011111010111110101","0000111010001110100011101000","0000110101001101010011010100","0000101011101010111010101110","0001000000000000000000000000","0000101011101010111010101110","0000001000010010000100100001","0000001100000011000000110000","0000100100001001000010010000","0000110101111101011111010111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111001101110011011100110","0000111101001111010011110100","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111011111110111111101111","0000111111111111111111111111","0000111010011110100111101001","0000110011101100111011001110","0000110001111100011111000111","0000110011001100110011001100","0000110111011101110111011101","0000111110001111100011111000","0000111010011110100111101001","0000100011001000110010001100","0000010011110100111101001111","0001000000000000000000000000","0000101101011011010110110101","0000101011101010111010101110","0000011010110110101101101011","0000100100001001000010010000","0000011101010111010101110101","0000001111010011110100111101","0000100000001000000010000000","0001000000000000000000000000","0000000000110000001100000011","0000010110000101100001011000","0000010110100101101001011010","0000110110101101101011011010","0000110010001100100011001000","0000110011111100111111001111","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111001111110011111100111","0000110110101101101011011010","0000101000101010001010100010","0000101010001010100010101000","0000101000011010000110100001","0000100110101001101010011010","0000110110101101101011011010","0000101101101011011010110110","0000100100111001001110010011","0000101111001011110010111100","0000101110101011101010111010","0000101010001010100010101000","0000110001011100010111000101","0000111010011110100111101001","0000110011111100111111001111","0000111100111111001111110011","0000101111001011110010111100","0000110010001100100011001000","0000101101101011011010110110","0000101100111011001110110011","0000100100111001001110010011","0000100011001000110010001100","0000010000100100001001000010","0000011110100111101001111010","0000000110000001100000011000","0000010101100101011001010110","0000011010000110100001101000","0000110000101100001011000010","0000111010011110100111101001","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000100101011001010110010101","0000101111001011110010111100","0000000101100001011000010110","0000000111110001111100011111","0000110111001101110011011100","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111110011111100111111001","0000111011111110111111101111","0000010011110100111101001111","0000010010000100100001001000","0000011111010111110101111101","0000110100001101000011010000","0000101011001010110010101100","0000111111111111111111111111","0000111101011111010111110101","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111110101111101011111010","0000101111111011111110111111","0000011101010111010101110101","0000100010111000101110001011","0000110110111101101111011011","0000110111011101110111011101","0000101011111010111110101111","0000011010100110101001101010","0000001010110010101100101011","0000010001100100011001000110","0000001010110010101100101011","0000000111110001111100011111","0000100101011001010110010101","0000111100011111000111110001","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111110001111100011111000","0000111111111111111111111111","0000111011001110110011101100","0000111011101110111011101110","0000010001000100010001000100","0000100011011000110110001101","0000110010001100100011001000","0000101100011011000110110001","0000110000101100001011000010","0000110111011101110111011101","0000111010001110100011101000","0000111001111110011111100111","0000100110101001101010011010","0000111010101110101011101010","0000011010110110101101101011","0000010010110100101101001011","0000010110010101100101011001","0000010001000100010001000100","0000100000001000000010000000","0000100000001000000010000000","0000100001101000011010000110","0000101010111010101110101011","0000100111111001111110011111","0000101010011010100110101001","0000101011001010110010101100","0000101010011010100110101001","0000100101011001010110010101","0000001011010010110100101101","0000011100110111001101110011","0000011101100111011001110110","0000100010101000101010001010","0000111000001110000011100000","0000111011011110110111101101","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111110011111100111111001","0000101110011011100110111001","0000011011110110111101101111","0000000010000000100000001000","0000101001001010010010100100","0000011000000110000001100000","0001000000000000000000000000","0000011010000110100001101000","0000101011011010110110101101","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111010011110100111101001","0000111101101111011011110110","0000111111111111111111111111","0000111011101110111011101110","0000111111001111110011111100","0000111010011110100111101001","0000111110111111101111111011","0000111100101111001011110010","0000111110101111101011111010","0000111101111111011111110111","0000110110011101100111011001","0000100110001001100010011000","0000110010011100100111001001","0000110111001101110011011100","0000100010001000100010001000","0000100100101001001010010010","0000010011100100111001001110","0000001011100010111000101110","0000100011011000110110001101","0000100110101001101010011010","0000100111111001111110011111","0000011110110111101101111011","0000001011010010110100101101","0000011110100111101001111010","0000000011110000111100001111","0000001010000010100000101000","0000010001010100010101000101","0000010010110100101101001011","0000110000001100000011000000","0000101001101010011010100110","0000111110111111101111111011","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111001011110010111100101","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111010001110100011101000","0000110110001101100011011000","0000100110001001100010011000","0000011110100111101001111010","0000010101000101010001010100","0000011101100111011001110110","0000100011011000110110001101","0000101010111010101110101011","0000100011101000111010001110","0000010101000101010001010100","0000011110100111101001111010","0000101100101011001010110010","0000101101111011011110110111","0000110000101100001011000010","0000101101001011010010110100","0000111001101110011011100110","0000110000001100000011000000","0000110010001100100011001000","0000100101101001011010010110","0000011111000111110001111100","0000100011101000111010001110","0000100010111000101110001011","0000010000110100001101000011","0000001011010010110100101101","0000001010110010101100101011","0000011011000110110001101100","0000011000100110001001100010","0000001100000011000000110000","0000100010111000101110001011","0000111101011111010111110101","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111101001111010011110100","0000101001011010010110100101","0000101010001010100010101000","0000001111010011110100111101","0000010011100100111001001110","0000110100101101001011010010","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000110000101100001011000010","0000000111110001111100011111","0000011010010110100101101001","0000100001101000011010000110","0000111011011110110111101101","0000110010111100101111001011","0000101101101011011010110110","0000111111111111111111111111","0000111011011110110111101101","0000111110001111100011111000","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000110111011101110111011101","0000100110001001100010011000","0000100101001001010010010100","0000100110101001101010011010","0000110010011100100111001001","0000110101101101011011010110","0000011110010111100101111001","0000011000000110000001100000","0000011000000110000001100000","0000010000010100000101000001","0000001110110011101100111011","0000001110000011100000111000","0000111011111110111111101111","0000111011111110111111101111","0000111111111111111111111111","0000111111011111110111111101","0000111000011110000111100001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000101001001010010010100100","0000010001010100010101000101","0000101010001010100010101000","0000100001111000011110000111","0000101001101010011010100110","0000101101101011011010110110","0000110101001101010011010100","0000111111111111111111111111","0000111001111110011111100111","0000101110011011100110111001","0000111011111110111111101111","0000110000101100001011000010","0000100100101001001010010010","0000101000001010000010100000","0000100001111000011110000111","0000011000110110001101100011","0000100010001000100010001000","0000100010001000100010001000","0000011010010110100101101001","0000011110010111100101111001","0000101010101010101010101010","0000101111011011110110111101","0000110001101100011011000110","0000100011101000111010001110","0000000010100000101000001010","0000010100100101001001010010","0000100100011001000110010001","0000110110111101101111011011","0000111001111110011111100111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000010100100101001001010010","0000010011110100111101001111","0000011001100110011001100110","0000110010011100100111001001","0000011001110110011101100111","0000000101000001010000010100","0000011110100111101001111010","0000110010011100100111001001","0000111101001111010011110100","0000111111011111110111111101","0000111100011111000111110001","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000110110101101101011011010","0000111101111111011111110111","0000110010101100101011001010","0000111011101110111011101110","0000111111111111111111111111","0000111110011111100111111001","0000111000001110000011100000","0000100011011000110110001101","0000110110111101101111011011","0000110101101101011011010110","0000100111111001111110011111","0000101100111011001110110011","0000011100100111001001110010","0000001011000010110000101100","0000010010100100101001001010","0000011001100110011001100110","0000101010101010101010101010","0000100010011000100110001001","0000001001000010010000100100","0000100100011001000110010001","0001000000000000000000000000","0000001001110010011100100111","0000010011100100111001001110","0000010000000100000001000000","0000011110010111100101111001","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111011001110110011101100","0000111101101111011011110110","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111011011110110111101101","0000110011101100111011001110","0000100010001000100010001000","0000010001110100011101000111","0000001110100011101000111010","0000010110010101100101011001","0000011011010110110101101101","0000011100000111000001110000","0000011010100110101001101010","0000011100110111001101110011","0000001101010011010100110101","0000010101100101011001010110","0000100110001001100010011000","0000110101111101011111010111","0000111100001111000011110000","0000110000101100001011000010","0000101100001011000010110000","0000100011001000110010001100","0000110000011100000111000001","0000101011111010111110101111","0000011110100111101001111010","0000010100110101001101010011","0000011000000110000001100000","0000011100000111000001110000","0000011001000110010001100100","0000001000000010000000100000","0000000011010000110100001101","0000001010110010101100101011","0000010001100100011001000110","0000010011000100110001001100","0000101110111011101110111011","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000100111111001111110011111","0000101100001011000010110000","0000001011000010110000101100","0000100001111000011110000111","0000110101111101011111010111","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000101011111010111110101111","0000000001000000010000000100","0000101110011011100110111001","0000110010011100100111001001","0000111011011110110111101101","0000111111111111111111111111","0000100111101001111010011110","0000111101101111011011110110","0000111100101111001011110010","0000111011011110110111101101","0000111111011111110111111101","0000111110111111101111111011","0000111011101110111011101110","0000111011111110111111101111","0000111000001110000011100000","0000101111101011111010111110","0000111000101110001011100010","0000101111011011110110111101","0000110010101100101011001010","0000110000111100001111000011","0000011110110111101101111011","0000010110110101101101011011","0000011010110110101101101011","0000010101010101010101010101","0000000000010000000100000001","0000100111001001110010011100","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111100111111001111110011","0000011111010111110101111101","0000001000110010001100100011","0000100001011000010110000101","0000010111110101111101011111","0000101101101011011010110110","0000101110011011100110111001","0000111010111110101111101011","0000111110001111100011111000","0000111011111110111111101111","0000110101001101010011010100","0000111011111110111111101111","0000111001001110010011100100","0000101110101011101010111010","0000111001101110011011100110","0000110011111100111111001111","0000101101101011011010110110","0000100101101001011010010110","0000101010111010101110101011","0000101101001011010010110100","0000101101001011010010110100","0000101101001011010010110100","0000101100101011001010110010","0000101101011011010110110101","0000010111010101110101011101","0000000011010000110100001101","0000010011100100111001001110","0000100010101000101010001010","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101111111011111110111","0000111001001110010011100100","0000000111010001110100011101","0000010100010101000101010001","0000001110000011100000111000","0000100110101001101010011010","0000110001111100011111000111","0000001101000011010000110100","0000001011110010111100101111","0000100000001000000010000000","0000110110011101100111011001","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000110000001100000011000000","0000111011011110110111101101","0000110000111100001111000011","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000101001011010010110100101","0000110010011100100111001001","0000101001101010011010100110","0000110000001100000011000000","0000100110011001100110011001","0000101100001011000010110000","0000011111000111110001111100","0001000000000000000000000000","0000011100100111001001110010","0000100100101001001010010010","0000011000000110000001100000","0000000011000000110000001100","0000010001010100010101000101","0000000011110000111100001111","0000001100100011001000110010","0000011111110111111101111111","0000011010000110100001101000","0000101011001010110010101100","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111100101111001011110010","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111001001110010011100100","0000100101111001011110010111","0000100010001000100010001000","0000010111110101111101011111","0000001100000011000000110000","0000000110000001100000011000","0000000000010000000100000001","0001000000000000000000000000","0001000000000000000000000000","0000000001110000011100000111","0000000000100000001000000010","0000001000010010000100100001","0000001110110011101100111011","0000010101010101010101010101","0000100000011000000110000001","0000100001111000011110000111","0000011001000110010001100100","0000010111010101110101011101","0000011010110110101101101011","0000011000100110001001100010","0000010100010101000101010001","0000011010000110100001101000","0000011011010110110101101101","0000010001000100010001000100","0000001010000010100000101000","0001000000000000000000000000","0000000010110000101100001011","0000001111010011110100111101","0000010101000101010001010100","0000010011110100111101001111","0000100101001001010010010100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000100110101001101010011010","0000110000101100001011000010","0000000000100000001000000010","0000100110101001101010011010","0000111100111111001111110011","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111100111111001111110011","0000111110011111100111111001","0000111110101111101011111010","0000011111010111110101111101","0000001100100011001000110010","0000110010111100101111001011","0000111001011110010111100101","0000111100111111001111110011","0000111111011111110111111101","0000111100001111000011110000","0000101111111011111110111111","0000111111101111111011111110","0000111111101111111011111110","0000111101011111010111110101","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110101001101010011010100","0000101111111011111110111111","0000111010011110100111101001","0000111100101111001011110010","0000110010011100100111001001","0000101011001010110010101100","0000100111111001111110011111","0000100010011000100110001001","0000011001000110010001100100","0000001111000011110000111100","0000000111100001111000011110","0000111100111111001111110011","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111000001110000011100000","0000010101100101011001010110","0000000011000000110000001100","0000011110000111100001111000","0000100100011001000110010001","0000101101011011010110110101","0000101001111010011110100111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111001101110011011100110","0000110111101101111011011110","0000111011101110111011101110","0000111110011111100111111001","0000101010001010100010101000","0000111101101111011011110110","0000111111011111110111111101","0000110010111100101111001011","0000110110011101100111011001","0000111100111111001111110011","0000111111011111110111111101","0000111100111111001111110011","0000111111001111110011111100","0000111111101111111011111110","0000011100100111001001110010","0000001010010010100100101001","0000010010100100101001001010","0000101001101010011010100110","0000111110001111100011111000","0000110111101101111011011110","0000111001111110011111100111","0000111101101111011011110110","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111011001110110011101100","0000110011011100110111001101","0000110001111100011111000111","0000100001111000011110000111","0000001011000010110000101100","0000011010010110100101101001","0000001011100010111000101110","0000010010100100101001001010","0000011100010111000101110001","0000100110001001100010011000","0000001001010010010100100101","0000001101100011011000110110","0000100011111000111110001111","0000111100011111000111110001","0000111111111111111111111111","0000111101111111011111110111","0000111011011110110111101101","0000111101111111011111110111","0000111110111111101111111011","0000111010111110101111101011","0000111001101110011011100110","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000110101001101010011010100","0000110011011100110111001101","0000111000001110000011100000","0000110101101101011011010110","0000111100101111001011110010","0000111110001111100011111000","0000111001001110010011100100","0000110001111100011111000111","0000110111101101111011011110","0000111101111111011111110111","0000101101101011011010110110","0000101010011010100110101001","0000101011101010111010101110","0000101010101010101010101010","0000010001100100011001000110","0001000000000000000000000000","0000010111110101111101011111","0000100010011000100110001001","0000000100110001001100010011","0000010011010100110101001101","0001000000000000000000000000","0000000100100001001000010010","0000010101110101011101010111","0000100011111000111110001111","0000110100101101001011010010","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111010101110101011101010","0000111111111111111111111111","0000111110001111100011111000","0000101011001010110010101100","0000100110101001101010011010","0000011110110111101101111011","0000001011000010110000101100","0000000010010000100100001001","0000000000110000001100000011","0000000110110001101100011011","0000010010110100101101001011","0000010101110101011101010111","0000011001110110011101100111","0000011011100110111001101110","0000001011010010110100101101","0000001100100011001000110010","0000001001100010011000100110","0000001100110011001100110011","0000000011000000110000001100","0001000000000000000000000000","0000001000110010001100100011","0000000110100001101000011010","0000001011110010111100101111","0000000100010001000100010001","0001000000000000000000000000","0001000000000000000000000000","0000000000110000001100000011","0000001001100010011000100110","0000001111000011110000111100","0000001000000010000000100000","0000000000010000000100000001","0000011100010111000101110001","0000101000011010000110100001","0000011100110111001101110011","0000111101011111010111110101","0000111101111111011111110111","0000111110101111101011111010","0000110111101101111011011110","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000100111011001110110011101","0000101001111010011110100111","0001000000000000000000000000","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111110111111101111111011","0000111100111111001111110011","0000110001101100011011000110","0000110111001101110011011100","0000111001011110010111100101","0000111100011111000111110001","0000001100000011000000110000","0000011111000111110001111100","0000100110111001101110011011","0000111110101111101011111010","0000111011111110111111101111","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111100101111001011110010","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111011111110111111101111","0000111010001110100011101000","0000101011001010110010101100","0000110000101100001011000010","0000111111111111111111111111","0000110111101101111011011110","0000111010101110101011101010","0000110000111100001111000011","0000111110111111101111111011","0000100100101001001010010010","0000101110101011101010111010","0000001011000010110000101100","0000010101010101010101010101","0000111100011111000111110001","0000111111111111111111111111","0000111010001110100011101000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000000001100000011000000110","0000001100110011001100110011","0000100001101000011010000110","0000101101101011011010110110","0000100010001000100010001000","0000101001111010011110100111","0000111101001111010011110100","0000111111111111111111111111","0000111001001110010011100100","0000111101101111011011110110","0000111000101110001011100010","0000111111101111111011111110","0000110110001101100011011000","0000110010111100101111001011","0000110011001100110011001100","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000011110100111101001111010","0000010010100100101001001010","0000001101000011010000110100","0000100100111001001110010011","0000111101001111010011110100","0000110110001101100011011000","0000101111001011110010111100","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111101011111010111110101","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110110011101100111011001","0000101010011010100110101001","0000100110101001101010011010","0001000000000000000000000000","0000010010000100100001001000","0000011101000111010001110100","0000100100101001001010010010","0000100000001000000010000000","0000100011111000111110001111","0000111111111111111111111111","0000111000011110000111100001","0000000100110001001100010011","0000001101100011011000110110","0000100111011001110110011101","0000111111001111110011111100","0000111111111111111111111111","0000111001101110011011100110","0000110101111101011111010111","0000110100011101000111010001","0000101011111010111110101111","0000110101101101011011010110","0000111101111111011111110111","0000111111111111111111111111","0000111101101111011011110110","0000111101011111010111110101","0000111110101111101011111010","0000101111101011111010111110","0000110001101100011011000110","0000110001011100010111000101","0000111110011111100111111001","0000111111111111111111111111","0000110001001100010011000100","0000110010001100100011001000","0000101110101011101010111010","0000111101101111011011110110","0000110110101101101011011010","0000101101101011011010110110","0000100100101001001010010010","0000110000101100001011000010","0000011110010111100101111001","0000000010010000100100001001","0000001101000011010000110100","0000001010000010100000101000","0000000000010000000100000001","0000001000010010000100100001","0001000000000000000000000000","0000001000110010001100100011","0000001010010010100100101001","0000011111010111110101111101","0000111111111111111111111111","0000111110101111101011111010","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000101100011011000110110001","0000100010011000100110001001","0000100111001001110010011100","0000011101110111011101110111","0000000010110000101100001011","0000000110000001100000011000","0000010111010101110101011101","0000011111110111111101111111","0000101000111010001110100011","0000011100100111001001110010","0000011011000110110001101100","0000011000010110000101100001","0000010100100101001001010010","0000100101101001011010010110","0000100101111001011110010111","0000010011100100111001001110","0000010001100100011001000110","0000010000110100001101000011","0000000011010000110100001101","0000000011000000110000001100","0000000010010000100100001001","0000001100110011001100110011","0000001111010011110100111101","0000010001110100011101000111","0000011010010110100101101001","0000100001111000011110000111","0000010101100101011001010110","0000011001010110010101100101","0000011101010111010101110101","0000111110011111100111111001","0000101100111011001110110011","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111101001111010011110100","0000111101111111011111110111","0000110110101101101011011010","0000100101011001010110010101","0000100000101000001010000010","0001000000000000000000000000","0000111001011110010111100101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111001111110011111100111","0000101100001011000010110000","0000110010011100100111001001","0000110100111101001111010011","0000101001011010010110100101","0000001101100011011000110110","0000100111111001111110011111","0000110101101101011011010110","0000111000001110000011100000","0000110101111101011111010111","0000111101111111011111110111","0000111011011110110111101101","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000110011111100111111001111","0000111001001110010011100100","0000011101100111011001110110","0000111001111110011111100111","0000110011101100111011001110","0000111111111111111111111111","0000110110111101101111011011","0000111110001111100011111000","0000111101101111011011110110","0000101111111011111110111111","0000101111101011111010111110","0000000001100000011000000110","0000100011011000110110001101","0000111100111111001111110011","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111110111111101111111011","0000000001000000010000000100","0000001010100010101000101010","0000100001101000011010000110","0000100101111001011110010111","0000100100011001000110010001","0000011001010110010101100101","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111010001110100011101000","0000111100111111001111110011","0000111101011111010111110101","0000110111101101111011011110","0000110001001100010011000100","0000110101101101011011010110","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111100011111000111110001","0000111110101111101011111010","0000111111111111111111111111","0000010010000100100001001000","0000001011000010110000101100","0000010010100100101001001010","0000011101110111011101110111","0000111100001111000011110000","0000111111001111110011111100","0000100111011001110110011101","0000111100101111001011110010","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000100001111000011110000111","0000101000001010000010100000","0000010010010100100101001001","0000000011110000111100001111","0000011010100110101001101010","0000111100011111000111110001","0000111000111110001111100011","0000101010001010100010101000","0000100100001001000010010000","0000110000011100000111000001","0000111010011110100111101001","0000110010101100101011001010","0000001101010011010100110101","0000001101100011011000110110","0000011110000111100001111000","0000011110000111100001111000","0000100101101001011010010110","0000100110011001100110011001","0000011110010111100101111001","0000110010001100100011001000","0000111001001110010011100100","0000111111001111110011111100","0000111110011111100111111001","0000111110011111100111111001","0000111000101110001011100010","0000111011011110110111101101","0000110010111100101111001011","0000110001011100010111000101","0000110110101101101011011010","0000111011101110111011101110","0000111111111111111111111111","0000101110001011100010111000","0000111000101110001011100010","0000100111001001110010011100","0000111010101110101011101010","0000111111111111111111111111","0000111010011110100111101001","0000100111001001110010011100","0000100010011000100110001001","0000101100011011000110110001","0000000110010001100100011001","0000000001010000010100000101","0000001100000011000000110000","0000000010100000101000001010","0000000010000000100000001000","0001000000000000000000000000","0000001101000011010000110100","0000001101100011011000110110","0000011111010111110101111101","0000111011111110111111101111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110011001100110011001100","0000011010000110100001101000","0000100011111000111110001111","0000100100111001001110010011","0001000000000000000000000000","0000011001110110011101100111","0000010010010100100101001001","0000011111000111110001111100","0000100101111001011110010111","0000011011010110110101101101","0000100000011000000110000001","0000011010100110101001101010","0000011011000110110001101100","0000011001110110011101100111","0000100010001000100010001000","0000100001011000010110000101","0000011000100110001001100010","0000011010100110101001101010","0000011100100111001001110010","0000010111000101110001011100","0000010000000100000001000000","0000010001010100010101000101","0000010100110101001101010011","0000010001000100010001000100","0000010111000101110001011100","0000010111110101111101011111","0000100011011000110110001101","0000100101011001010110010101","0000011000110110001101100011","0000110000101100001011000010","0000110110111101101111011011","0000111101001111010011110100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111110001111100011111000","0000101111011011110110111101","0000100011011000110110001101","0000010110010101100101011001","0001000000000000000000000000","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111100001111000011110000","0000110111101101111011011110","0000100000111000001110000011","0000100000101000001010000010","0000110001011100010111000101","0000010001100100011001000110","0000011010000110100001101000","0000100011111000111110001111","0000100101111001011110010111","0000110001011100010111000101","0000111111001111110011111100","0000111110011111100111111001","0000111110011111100111111001","0000111111101111111011111110","0000111110011111100111111001","0000111101011111010111110101","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000110000011100000111000001","0000111001001110010011100100","0000101111001011110010111100","0000111011101110111011101110","0000111000111110001111100011","0000111010001110100011101000","0000111011001110110011101100","0000111111011111110111111101","0000111111111111111111111111","0000110011101100111011001110","0000101001011010010110100101","0001000000000000000000000000","0000110011101100111011001110","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111101001111010011110100","0001000000000000000000000000","0001000000000000000000000000","0000011000010110000101100001","0000100011101000111010001110","0000100111101001111010011110","0000010010110100101101001011","0000111110111111101111111011","0000111111111111111111111111","0000111011111110111111101111","0000110011001100110011001100","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111111101111111011111110","0000111100011111000111110001","0000110111011101110111011101","0000110110011101100111011001","0000111010111110101111101011","0000111111111111111111111111","0000111100011111000111110001","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000011110000111100001111000","0000001000010010000100100001","0000000111100001111000011110","0000100001001000010010000100","0000111111111111111111111111","0000110100101101001011010010","0000110110101101101011011010","0000110001011100010111000101","0000111111111111111111111111","0000111011011110110111101101","0000111110101111101011111010","0000111111111111111111111111","0000111011001110110011101100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000101111101011111010111110","0000011001000110010001100100","0000010001100100011001000110","0000000110110001101100011011","0000011101000111010001110100","0000110001101100011011000110","0000111111111111111111111111","0000111111111111111111111111","0000101111001011110010111100","0000101101011011010110110101","0000101111001011110010111100","0000111110101111101011111010","0000110010011100100111001001","0000110001001100010011000100","0000010101100101011001010110","0000001001100010011000100110","0000010010000100100001001000","0000010110100101101001011010","0000101111101011111010111110","0000110110001101100011011000","0000111111001111110011111100","0000111111101111111011111110","0000111010101110101011101010","0000111101001111010011110100","0000111010011110100111101001","0000110011101100111011001110","0000110110001101100011011000","0000101000111010001110100011","0000101110001011100010111000","0000101011011010110110101101","0000110010011100100111001001","0000111111111111111111111111","0000101101101011011010110110","0000110110101101101011011010","0000101001001010010010100100","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110001001100010011000100","0000100010011000100110001001","0000100111011001110110011101","0000010010110100101101001011","0000000110010001100100011001","0000001011000010110000101100","0000000100000001000000010000","0000010010010100100101001001","0001000000000000000000000000","0000001000000010000000100000","0000000111010001110100011101","0000100000001000000010000000","0000111111011111110111111101","0000111110001111100011111000","0000111111001111110011111100","0000111110101111101011111010","0000111101001111010011110100","0000101000011010000110100001","0000101110001011100010111000","0000100001101000011010000110","0000101001011010010110100101","0000011110000111100001111000","0000101110111011101110111011","0000101000011010000110100001","0000101100011011000110110001","0000110100101101001011010010","0000101111101011111010111110","0000111100001111000011110000","0000101110111011101110111011","0000101010001010100010101000","0000111100011111000111110001","0000111111001111110011111100","0000111001101110011011100110","0000110111001101110011011100","0000101010101010101010101010","0000100000011000000110000001","0000100000111000001110000011","0000010000010100000101000001","0000010001010100010101000101","0000010001010100010101000101","0000001101100011011000110110","0000010000010100000101000001","0000010110010101100101011001","0000101110001011100010111000","0000101101011011010110110101","0000101000101010001010100010","0000111000111110001111100011","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111111011111110111111101","0000111111001111110011111100","0000111110001111100011111000","0000111110111111101111111011","0000111101011111010111110101","0000101100001011000010110000","0000100011111000111110001111","0000001001000010010000100100","0000010110100101101001011010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000110111011101110111011101","0000101010101010101010101010","0000010110110101101101011011","0000011100010111000101110001","0000011000110110001101100011","0000010010010100100101001001","0000011111010111110101111101","0000011111100111111001111110","0000100011111000111110001111","0000110101101101011011010110","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111001011110010111100101","0000110010101100101011001010","0000111001101110011011100110","0000110101101101011011010110","0000110010111100101111001011","0000101010101010101010101010","0000110000101100001011000010","0000111010001110100011101000","0000110110101101101011011010","0000111111111111111111111111","0000111100001111000011110000","0000111001011110010111100101","0000111110001111100011111000","0000110101111101011111010111","0000010000010100000101000001","0000001100010011000100110001","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0001000000000000000000000000","0000001000110010001100100011","0000001001110010011100100111","0000101010111010101110101011","0000011111000111110001111100","0000100011101000111010001110","0000110110011101100111011001","0000111111011111110111111101","0000111111111111111111111111","0000100110111001101110011011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111100001111000011110000","0000111111111111111111111111","0000111110011111100111111001","0000111110111111101111111011","0000111111001111110011111100","0000100010011000100110001001","0000000111100001111000011110","0000000010010000100100001001","0000010011110100111101001111","0000100110111001101110011011","0000111000101110001011100010","0000110101111101011111010111","0000100111001001110010011100","0000111011101110111011101110","0000111110001111100011111000","0000111111111111111111111111","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111000011110000111100001","0000011110000111100001111000","0000010001010100010101000101","0000000110010001100100011001","0000001110100011101000111010","0000100010011000100110001001","0000110111101101111011011110","0000111110101111101011111010","0000111111111111111111111111","0000110111111101111111011111","0000110100011101000111010001","0000101001101010011010100110","0000111100001111000011110000","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000101101101011011010110110","0000011011000110110001101100","0000011110100111101001111010","0000010010110100101101001011","0000100011001000110010001100","0000100110111001101110011011","0000101101011011010110110101","0000110010011100100111001001","0000111101101111011011110110","0000111111001111110011111100","0000110000011100000111000001","0000110000101100001011000010","0000100001011000010110000101","0000011111010111110101111101","0000011101010111010101110101","0000110010011100100111001001","0000110010011100100111001001","0000101101001011010010110100","0000110101001101010011010100","0000110100101101001011010010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111011011110110111101101","0000101011101010111010101110","0000011111110111111101111111","0000011110100111101001111010","0000001001000010010000100100","0000001111010011110100111101","0000000000010000000100000001","0000010001100100011001000110","0000000011010000110100001101","0000000110010001100100011001","0000001110000011100000111000","0000100101101001011010010110","0000111100011111000111110001","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000110000011100000111000001","0000110011011100110111001101","0000101110101011101010111010","0000101110111011101110111011","0000101100001011000010110000","0000111011001110110011101100","0000110001001100010011000100","0000110100001101000011010000","0000110101001101010011010100","0000111010111110101111101011","0000110100111101001111010011","0000111111111111111111111111","0000110101001101010011010100","0000110100111101001111010011","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111000001110000011100000","0000101100101011001010110010","0000101001011010010110100101","0000011101100111011001110110","0000011000100110001001100010","0000100001101000011010000110","0000101010111010101110101011","0000101001101010011010100110","0000101001011010010110100101","0000111010011110100111101001","0000110001001100010011000100","0000110100011101000111010001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111110111111101111111011","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111001001110010011100100","0000100110001001100010011000","0000100101111001011110010111","0000000010110000101100001011","0000011111000111110001111100","0000111100111111001111110011","0000111111101111111011111110","0000111000111110001111100011","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000011100000111000001110000","0000010000010100000101000001","0000010001100100011001000110","0000000011110000111100001111","0000011101010111010101110101","0000011101100111011001110110","0000011000000110000001100000","0000101000111010001110100011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111100011111000111110001","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000110010011100100111001001","0000110011001100110011001100","0000101111111011111110111111","0000110100001101000011010000","0000110011111100111111001111","0000111100101111001011110010","0000111100001111000011110000","0000111000101110001011100010","0000110000011100000111000001","0000111101111111011111110111","0000111010011110100111101001","0000111011011110110111101101","0000101001011010010110100101","0000010001100100011001000110","0000100111011001110110011101","0000111111101111111011111110","0000111110001111100011111000","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111100111111001111110011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000101010101010101010101010","0000000010100000101000001010","0000001000100010001000100010","0001000000000000000000000000","0000011101010111010101110101","0000011100100111001001110010","0000100010111000101110001011","0000100110001001100010011000","0000111110101111101011111010","0000111110111111101111111011","0000101000011010000110100001","0000110111111101111111011111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111011101110111011101110","0000111100011111000111110001","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000101111011011110110111101","0000001101000011010000110100","0001000000000000000000000000","0000001001000010010000100100","0000100000001000000010000000","0000100010001000100010001000","0000101000001010000010100000","0000110100001101000011010000","0000101100101011001010110010","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000110001101100011011000110","0000011100100111001001110010","0000010011010100110101001101","0000001010000010100000101000","0000011100110111001101110011","0000101011101010111010101110","0000111110001111100011111000","0000111111001111110011111100","0000111101111111011111110111","0000111101111111011111110111","0000110101101101011011010110","0000101001001010010010100100","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000111100111111001111110011","0000111101101111011011110110","0000110011101100111011001110","0000100001101000011010000110","0000110011011100110111001101","0000110001001100010011000100","0000110100001101000011010000","0000111010011110100111101001","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000101100101011001010110010","0000101100101011001010110010","0000101010111010101110101011","0000011100010111000101110001","0000010001000100010001000100","0000010000110100001101000011","0000101101101011011010110110","0000011111110111111101111111","0000111010111110101111101011","0000101110111011101110111011","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000011101100111011001110110","0000100001001000010010000100","0000001010010010100100101001","0000010110000101100001011000","0001000000000000000000000000","0000001011010010110100101101","0000000001100000011000000110","0000001001010010010100100101","0000011100000111000001110000","0000100001111000011110000111","0000110111011101110111011101","0000111111111111111111111111","0000111110011111100111111001","0000111110111111101111111011","0000111000001110000011100000","0000111011001110110011101100","0000101101101011011010110110","0000110010111100101111001011","0000111010001110100011101000","0000111100011111000111110001","0000110000101100001011000010","0000111000111110001111100011","0000111011101110111011101110","0000111101001111010011110100","0000111000101110001011100010","0000111110111111101111111011","0000110110101101101011011010","0000111101101111011011110110","0000111100101111001011110010","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111011001110110011101100","0000100100111001001110010011","0000100110001001100010011000","0000100000101000001010000010","0000100111101001111010011110","0000110001111100011111000111","0000110010001100100011001000","0000111000011110000111100001","0000111111111111111111111111","0000110111001101110011011100","0000111011111110111111101111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110001001100010011000100","0000100110001001100010011000","0000100000111000001110000011","0001000000000000000000000000","0000100101001001010010010100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000001011000010110000101100","0000010001010100010101000101","0001000000000000000000000000","0000010001110100011101000111","0000100010101000101010001010","0000011011010110110101101101","0000100100011001000110010001","0000111011001110110011101100","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111001011110010111100101","0000101100001011000010110000","0000011110010111100101111001","0000100101101001011010010110","0000101000001010000010100000","0000100111011001110110011101","0000110010001100100011001000","0000111111011111110111111101","0000101110001011100010111000","0000111010101110101011101010","0000111001001110010011100100","0000110101011101010111010101","0000111111111111111111111111","0000110001011100010111000101","0000101001111010011110100111","0000001011100010111000101110","0000111011101110111011101110","0000111111001111110011111100","0000111100011111000111110001","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101011111010111110101","0000111111111111111111111111","0000011101100111011001110110","0000100011001000110010001100","0000001001010010010100100101","0000000011110000111100001111","0000010100010101000101010001","0000011101110111011101110111","0000010110110101101101011011","0000000111000001110000011100","0000101101011011010110110101","0000101111101011111010111110","0000010111110101111101011111","0000101001011010010110100101","0000110011001100110011001100","0000101101101011011010110110","0000101100111011001110110011","0000110011011100110111001101","0000111001101110011011100110","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000010101010101010101010101","0000000000100000001000000010","0000010001000100010001000100","0000000110010001100100011001","0000010000100100001001000010","0000001110010011100100111001","0000100000111000001110000011","0000100101001001010010010100","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000101011101010111010101110","0000011001010110010101100101","0000001110100011101000111010","0000000111110001111100011111","0000011010110110101101101011","0000101011011010110110101101","0000111110111111101111111011","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111001101110011011100110","0000101011011010110110101101","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000110100001101000011010000","0000111101111111011111110111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000110001011100010111000101","0000011110010111100101111001","0000100100111001001110010011","0000011101000111010001110100","0000001000010010000100100001","0000011000010110000101100001","0000011111000111110001111100","0000101111011011110110111101","0000101110011011100110111001","0000111011011110110111101101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000100101101001011010010110","0000011111110111111101111111","0000010000110100001101000011","0000010100000101000001010000","0000000001010000010100000101","0000001101000011010000110100","0000000000010000000100000001","0000001101010011010100110101","0000011101110111011101110111","0000011111000111110001111100","0000110011001100110011001100","0000111100111111001111110011","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111100011111000111110001","0000101101101011011010110110","0000110001111100011111000111","0000111111111111111111111111","0000110110001101100011011000","0000111001011110010111100101","0000111011001110110011101100","0000111100101111001011110010","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000100000101000001010000010","0000100000011000000110000001","0000011111000111110001111100","0000100110011001100110011001","0000101111111011111110111111","0000110011111100111111001111","0000111101011111010111110101","0000111010001110100011101000","0000111011111110111111101111","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111111011111110111111101","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000110101111101011111010111","0000101010001010100010101000","0000100101011001010110010101","0000001111100011111000111110","0000000001100000011000000110","0000111001111110011111100111","0000111111001111110011111100","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000101011101010111010101110","0000000111100001111000011110","0000010011100100111001001110","0000000111110001111100011111","0000010011010100110101001101","0000100110001001100010011000","0000100101001001010010010100","0000110101111101011111010111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111011111110111111101111","0000110101101101011011010110","0000010101110101011101010111","0000100000101000001010000010","0000001011000010110000101100","0000001000000010000000100000","0000011001100110011001100110","0000100110001001100010011000","0000100100011001000110010001","0000101011011010110110101101","0000110001111100011111000111","0000111100101111001011110010","0000110100111101001111010011","0000110011111100111111001111","0000110000111100001111000011","0000001110010011100100111001","0000101010011010100110101001","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101001111010011110100","0000111110011111100111111001","0001000000000000000000000000","0000010110010101100101011001","0000000101100001011000010110","0001000000000000000000000000","0000010100100101001001010010","0000010100000101000001010000","0000010110000101100001011000","0000011011100110111001101110","0000011001110110011101100111","0000110111001101110011011100","0000010100010101000101010001","0000011100110111001101110011","0000110001101100011011000110","0000101111011011110110111101","0000101011101010111010101110","0000101000001010000010100000","0000100110111001101110011011","0000101001011010010110100101","0000101110011011100110111001","0000110010011100100111001001","0000111000111110001111100011","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111011101110111011101110","0000100100101001001010010010","0000001101010011010100110101","0000000111010001110100011101","0000011011010110110101101101","0000010010000100100001001000","0000000101000001010000010100","0000001100110011001100110011","0000010011000100110001001100","0000011011110110111101101111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000101100101011001010110010","0000011100110111001101110011","0000001111110011111100111111","0000010001000100010001000100","0000011110000111100001111000","0000100110101001101010011010","0000111010111110101111101011","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000101100111011001110110011","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111000111110001111100011","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111010011110100111101001","0000111101101111011011110110","0000111111011111110111111101","0000111111001111110011111100","0000011010100110101001101010","0000011110000111100001111000","0000010110110101101101011011","0000001000010010000100100001","0000010100010101000101010001","0000010000100100001001000010","0000101000011010000110100001","0000100011011000110110001101","0000111101011111010111110101","0000111100011111000111110001","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111100001111000011110000","0000110011001100110011001100","0000100001111000011110000111","0000011010110110101101101011","0000001010010010100100101001","0001000000000000000000000000","0000000101000001010000010100","0000001010100010101000101010","0000010011010100110101001101","0000010111010101110101011101","0000101111101011111010111110","0000101000101010001010100010","0000110111011101110111011101","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000101101011011010110110101","0000110110101101101011011010","0000111111111111111111111111","0000111010001110100011101000","0000111100101111001011110010","0000111010111110101111101011","0000111100001111000011110000","0000111011111110111111101111","0000111111111111111111111111","0000111101111111011111110111","0000111011011110110111101101","0000111111011111110111111101","0000111101111111011111110111","0000111100111111001111110011","0000111011101110111011101110","0000111111111111111111111111","0000111100101111001011110010","0000111011101110111011101110","0000100111001001110010011100","0000011110100111101001111010","0000011111110111111101111111","0000101110001011100010111000","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111111101111111011111110","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111011011110110111101101","0000101100111011001110110011","0000100101001001010010010100","0000010111010101110101011101","0000000001010000010100000101","0000100000011000000110000001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111101101111011011110110","0000100111111001111110011111","0000010111010101110101011101","0000000011000000110000001100","0000001100000011000000110000","0000011100110111001101110011","0000101000101010001010100010","0000110110011101100111011001","0000111111101111111011111110","0000111010011110100111101001","0000111110001111100011111000","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000110100101101001011010010","0000011111010111110101111101","0000001110110011101100111011","0000000110100001101000011010","0000000111010001110100011101","0001000000000000000000000000","0001000000000000000000000000","0000000010000000100000001000","0001000000000000000000000000","0000010101010101010101010101","0000010011110100111101001111","0000001100000011000000110000","0000100010011000100110001001","0000110100011101000111010001","0000101100101011001010110010","0000111100001111000011110000","0000101001111010011110100111","0000011110000111100001111000","0000001111000011110000111100","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111011111110111111101","0000101010101010101010101010","0001000000000000000000000000","0001000000000000000000000000","0000001110000011100000111000","0000001110110011101100111011","0000100010001000100010001000","0000101001001010010010100100","0000011100000111000001110000","0000000011110000111100001111","0000011010000110100001101000","0000010101010101010101010101","0000001000100010001000100010","0000010010000100100001001000","0000011011100110111001101110","0000011011000110110001101100","0000010101100101011001010110","0000010010010100100101001001","0000011100000111000001110000","0000101101001011010010110100","0000110100101101001011010010","0000110001111100011111000111","0000110011111100111111001111","0000110010111100101111001011","0000111010011110100111101001","0000111111111111111111111111","0000111110111111101111111011","0000110110011101100111011001","0000011111000111110001111100","0000000011110000111100001111","0000011101000111010001110100","0000101110101011101010111010","0000101110111011101110111011","0000011000110110001101100011","0000010101100101011001010110","0000011001000110010001100100","0000011111010111110101111101","0000100110001001100010011000","0000101011101010111010101110","0000110010101100101011001010","0000101101101011011010110110","0000100111101001111010011110","0000100000111000001110000011","0000001000110010001100100011","0000010111100101111001011110","0000011001000110010001100100","0000110101001101010011010100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111101111111011111110111","0000110011111100111111001111","0000111101111111011111110111","0000111101011111010111110101","0000111111001111110011111100","0000111010011110100111101001","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111010101110101011101010","0000110100111101001111010011","0000001111110011111100111111","0000000111100001111000011110","0000100001111000011110000111","0000001100000011000000110000","0000000011010000110100001101","0000001111000011110000111100","0000100110101001101010011010","0000100001001000010010000100","0000111010111110101111101011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111100001111000011110000","0000111011101110111011101110","0000100110101001101010011010","0000011110110111101101111011","0000000101000001010000010100","0000000100000001000000010000","0001000000000000000000000000","0000001111110011111100111111","0000011101100111011001110110","0000011000000110000001100000","0000110101011101010111010101","0000100001101000011010000110","0000110100001101000011010000","0000111110111111101111111011","0000111111011111110111111101","0000111111011111110111111101","0000111101111111011111110111","0000111001111110011111100111","0000110110011101100111011001","0000111110111111101111111011","0000111101101111011011110110","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111101011111010111110101","0000111010011110100111101001","0000100101011001010110010101","0000100101101001011010010110","0000100110111001101110011011","0000110010011100100111001001","0000110100111101001111010011","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111010101110101011101010","0000101010001010100010101000","0000011111100111111001111110","0000001010110010101100101011","0000000101110001011100010111","0000111100101111001011110010","0000111011101110111011101110","0000111111111111111111111111","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000110010011100100111001001","0000101011111010111110101111","0000010001100100011001000110","0000001100000011000000110000","0000011000110110001101100011","0000100111011001110110011101","0000100110101001101010011010","0000111111001111110011111100","0000111111111111111111111111","0000111011101110111011101110","0000111100111111001111110011","0000111110111111101111111011","0000111100011111000111110001","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000110110101101101011011010","0000101000011010000110100001","0000011100010111000101110001","0000001110100011101000111010","0000001101000011010000110100","0000000100000001000000010000","0000000100110001001100010011","0000001000110010001100100011","0000001010000010100000101000","0000010000010100000101000001","0000001100100011001000110010","0000000100110001001100010011","0000001011110010111100101111","0000010000000100000001000000","0000001001010010010100100101","0000011100100111001001110010","0000111000001110000011100000","0000111000111110001111100011","0000100011001000110010001100","0000100100011001000110010001","0000000000100000001000000010","0000110000011100000111000001","0000111111111111111111111111","0000111111101111111011111110","0000111100101111001011110010","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011111110111111101111","0000001100010011000100110001","0000100110001001100010011000","0000001010110010101100101011","0000000001000000010000000100","0000000101000001010000010100","0000011111110111111101111111","0000011111100111111001111110","0000100010011000100110001001","0000010101010101010101010101","0000001100010011000100110001","0000100011001000110010001100","0000001100100011001000110010","0000010100100101001001010010","0000101100111011001110110011","0000110100111101001111010011","0000111010111110101111101011","0000111001101110011011100110","0000110110101101101011011010","0000110101101101011011010110","0000110100111101001111010011","0000110011001100110011001100","0000110111011101110111011101","0000101110101011101010111010","0000101110001011100010111000","0000111111011111110111111101","0000111111111111111111111111","0000111011101110111011101110","0000101100101011001010110010","0000100111101001111010011110","0000000000110000001100000011","0000100111111001111110011111","0000100111111001111110011111","0000110010101100101011001010","0000010111100101111001011110","0000010100010101000101010001","0000010111100101111001011110","0000110100111101001111010011","0000111011001110110011101100","0000111110001111100011111000","0000110101111101011111010111","0000100101101001011010010110","0000100011011000110110001101","0001000000000000000000000000","0000011011100110111001101110","0000010101010101010101010101","0000110100111101001111010011","0000111010101110101011101010","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111100101111001011110010","0000111101011111010111110101","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111101001111010011110100","0000111111101111111011111110","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000101101001011010010110100","0000100010001000100010001000","0000011011010110110101101101","0000010101000101010001010100","0000010000100100001001000010","0000001111010011110100111101","0000001111000011110000111100","0000010010000100100001001000","0000010111110101111101011111","0000101011011010110110101101","0000011011110110111101101111","0000111010011110100111101001","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000101001111010011110100111","0000011100100111001001110010","0000000110100001101000011010","0000010000110100001101000011","0000000101000001010000010100","0000000110100001101000011010","0000100110111001101110011011","0000011101110111011101110111","0000100010101000101010001010","0000100101001001010010010100","0000110001001100010011000100","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000111111011111110111111101","0000111100101111001011110010","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111110101111101011111010","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111110101111101011111010","0000111100001111000011110000","0000111000011110000111100001","0000010111100101111001011110","0000101011011010110110101101","0000100111111001111110011111","0000110111111101111111011111","0000111000011110000111100001","0000111111111111111111111111","0000110001011100010111000101","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000101010111010101110101011","0000011010000110100001101000","0000001100000011000000110000","0000010010110100101101001011","0000111100101111001011110010","0000111111111111111111111111","0000111101011111010111110101","0000111011111110111111101111","0000111101011111010111110101","0000111101011111010111110101","0000110101001101010011010100","0000101010001010100010101000","0000100000111000001110000011","0000011000100110001001100010","0000100111111001111110011111","0000100110001001100010011000","0000101100001011000010110000","0000111011001110110011101100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111000101110001011100010","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000101011101010111010101110","0000010011110100111101001111","0000001001000010010000100100","0000000010100000101000001010","0000001100100011001000110010","0000100110101001101010011010","0000100101001001010010010100","0000001101010011010100110101","0000010111100101111001011110","0000011100010111000101110001","0000001010010010100100101001","0000010111110101111101011111","0000001100110011001100110011","0000010000000100000001000000","0000001010100010101000101010","0000010001010100010101000101","0000100101101001011010010110","0000101110101011101010111010","0000110001001100010011000100","0000100110001001100010011000","0000001101100011011000110110","0000100011001000110010001100","0000111101011111010111110101","0000111111011111110111111101","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101111111011111110111","0000100101001001010010010100","0000000001000000010000000100","0000100101001001010010010100","0000010101010101010101010101","0000101110001011100010111000","0000011011010110110101101101","0000010101010101010101010101","0000000110110001101100011011","0000001011110010111100101111","0000001000100010001000100010","0000001001100010011000100110","0000001111010011110100111101","0000000110110001101100011011","0000001101010011010100110101","0000010000110100001101000011","0000011011000110110001101100","0000011011000110110001101100","0000101110101011101010111010","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111000011110000111100001","0000111011011110110111101101","0000011110010111100101111001","0000111000101110001011100010","0000111111111111111111111111","0000111111001111110011111100","0000111010111110101111101011","0000110111001101110011011100","0000110001001100010011000100","0000010101000101010001010100","0000011100010111000101110001","0000110101011101010111010101","0000101000001010000010100000","0000011111010111110101111101","0000011010010110100101101001","0000110100011101000111010001","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000100101111001011110010111","0000101001101010011010100110","0001000000000000000000000000","0000011010100110101001101010","0000011000110110001101100011","0000101110111011101110111011","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111010101110101011101010","0000111011101110111011101110","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111000001110000011100000","0000101110011011100110111001","0000100101011001010110010101","0000100010101000101010001010","0000100000101000001010000010","0000011001000110010001100100","0000001110110011101100111011","0000000111110001111100011111","0000011010000110100001101000","0000011011110110111101101111","0000010100100101001001010010","0000010101110101011101010111","0000101010111010101110101011","0000011011000110110001101100","0000111101111111011111110111","0000111100101111001011110010","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000100100011001000110010001","0000011001110110011101100111","0000010000000100000001000000","0000010000000100000001000000","0001000000000000000000000000","0000000111110001111100011111","0000110001101100011011000110","0000011110100111101001111010","0000100110101001101010011010","0000110010101100101011001010","0000100111111001111110011111","0000111001101110011011100110","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111101101111011011110110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111010101110101011101010","0000111010111110101111101011","0000011001100110011001100110","0000011110110111101101111011","0000100111001001110010011100","0000110010011100100111001001","0000111101111111011111110111","0000111110011111100111111001","0000111000111110001111100011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111100011111000111110001","0000111101011111010111110101","0000111111111111111111111111","0000111110001111100011111000","0000111010101110101011101010","0000111000111110001111100011","0000100100011001000110010001","0000011101010111010101110101","0000000110100001101000011010","0000101000111010001110100011","0000111101011111010111110101","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000110110101101101011011010","0000100111001001110010011100","0000101010111010101110101011","0000101111011011110110111101","0000101111111011111110111111","0000100100011001000110010001","0000110101001101010011010100","0000101111101011111010111110","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111100011111000111110001","0000111110011111100111111001","0000111110001111100011111000","0000111101101111011011110110","0000110011001100110011001100","0000011011000110110001101100","0000011001000110010001100100","0000010000000100000001000000","0000010000100100001001000010","0000111100001111000011110000","0000111100001111000011110000","0000011101110111011101110111","0000011000000110000001100000","0000010010100100101001001010","0000100001001000010010000100","0000011010100110101001101010","0000011011100110111001101110","0000100110001001100010011000","0000000011100000111000001110","0000001110010011100100111001","0000010011110100111101001111","0000011010010110100101101001","0000101100011011000110110001","0000111110001111100011111000","0000011010110110101101101011","0000011010110110101101101011","0000001000100010001000100010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000110111111101111111011111","0000000000100000001000000010","0000101111111011111110111111","0000100001101000011010000110","0000111000001110000011100000","0000110100111101001111010011","0000110011011100110111001101","0000100111111001111110011111","0000101110001011100010111000","0000100001011000010110000101","0000100000011000000110000001","0000100011001000110010001100","0000110101111101011111010111","0000011101000111010001110100","0000011100100111001001110010","0000110101011101010111010101","0000111011001110110011101100","0000110001101100011011000110","0000110001111100011111000111","0000100111001001110010011100","0000111100011111000111110001","0000111111111111111111111111","0000111001011110010111100101","0000111110101111101011111010","0000111001101110011011100110","0000111100111111001111110011","0000101011001010110010101100","0000111100001111000011110000","0000111111101111111011111110","0000111111111111111111111111","0000110101001101010011010100","0000111011101110111011101110","0000110011111100111111001111","0000010100110101001101010011","0000011101110111011101110111","0000110110011101100111011001","0000100001101000011010000110","0000100101001001010010010100","0000110100111101001111010011","0000111111011111110111111101","0000111111111111111111111111","0000111101111111011111110111","0000101001001010010010100100","0000100000001000000010000000","0000001001100010011000100110","0000011111010111110101111101","0000011001100110011001100110","0000100010101000101010001010","0000110100101101001011010010","0000111101001111010011110100","0000111000001110000011100000","0000111111111111111111111111","0000111011111110111111101111","0000111100001111000011110000","0000101111111011111110111111","0000110001101100011011000110","0000110101101101011011010110","0000111110101111101011111010","0000111101111111011111110111","0000111000101110001011100010","0000101010101010101010101010","0000100111011001110110011101","0000100111011001110110011101","0000010111000101110001011100","0000100101101001011010010110","0000100110001001100010011000","0000010011000100110001001100","0000000111010001110100011101","0000001101100011011000110110","0000010011100100111001001110","0000010001000100010001000100","0000100110011001100110011001","0000001011010010110100101101","0000011011000110110001101100","0000010001100100011001000110","0000110101101101011011010110","0000011100000111000001110000","0000111001011110010111100101","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111110111111101111111011","0000111101111111011111110111","0000110001001100010011000100","0000100101011001010110010101","0000100011001000110010001100","0000011100100111001001110010","0000010001100100011001000110","0000000001110000011100000111","0000000111010001110100011101","0000101001001010010010100100","0000011011000110110001101100","0000100001011000010110000101","0000111010001110100011101000","0000111011001110110011101100","0000111000001110000011100000","0000111011101110111011101110","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111011111110111111101111","0000111101111111011111110111","0000110111001101110011011100","0000101010111010101110101011","0000100100111001001110010011","0000011001100110011001100110","0000101110111011101110111011","0000100111001001110010011100","0000110100001101000011010000","0000110110001101100011011000","0000110011001100110011001100","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110000101100001011000010","0000100111111001111110011111","0000010100110101001101010011","0000010001000100010001000100","0000100110101001101010011010","0000111001011110010111100101","0000111000101110001011100010","0000111110101111101011111010","0000111101101111011011110110","0000111101101111011011110110","0000111110001111100011111000","0000111001001110010011100100","0000101110111011101110111011","0000110010011100100111001001","0000111010001110100011101000","0000111011111110111111101111","0000110011111100111111001111","0000110010001100100011001000","0000110110111101101111011011","0000111100011111000111110001","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111011111110111111101","0000111111111111111111111111","0000110100101101001011010010","0000101010101010101010101010","0000011000110110001101100011","0000010111000101110001011100","0000000101110001011100010111","0000111001001110010011100100","0000111011011110110111101101","0000111111001111110011111100","0000101000111010001110100011","0000011010010110100101101001","0000011001110110011101100111","0000010101010101010101010101","0000011110110111101101111011","0000011111100111111001111110","0000111010011110100111101001","0000010111110101111101011111","0000000001110000011100000111","0000001101100011011000110110","0000011100000111000001110000","0000100000111000001110000011","0000111111111111111111111111","0000100010111000101110001011","0000011011100110111001101110","0000000000100000001000000010","0000110001111100011111000111","0000111100101111001011110010","0000111110101111101011111010","0000111110011111100111111001","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000010010100100101001001010","0000010100100101001001010010","0000111100011111000111110001","0000101100101011001010110010","0000111111011111110111111101","0000111101011111010111110101","0000110111001101110011011100","0000110010111100101111001011","0000100100001001000010010000","0000100011111000111110001111","0000011000010110000101100001","0000011000010110000101100001","0000110100101101001011010010","0000100000101000001010000010","0000011001110110011101100111","0000110011011100110111001101","0000111110011111100111111001","0000110000111100001111000011","0000111111111111111111111111","0000111001011110010111100101","0000111011011110110111101101","0000111110111111101111111011","0000111110111111101111111011","0000111101001111010011110100","0000111111111111111111111111","0000111110011111100111111001","0000101110111011101110111011","0000111000011110000111100001","0000111100101111001011110010","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111010111110101111101011","0000101010001010100010101000","0000100011011000110110001101","0000100111101001111010011110","0000101011101010111010101110","0000100111011001110110011101","0000110010101100101011001010","0000111100001111000011110000","0000111101001111010011110100","0000111111111111111111111111","0000110110011101100111011001","0000011000100110001001100010","0000011000010110000101100001","0000100011101000111010001110","0000100001111000011110000111","0000011000000110000001100000","0000100010111000101110001011","0000110101001101010011010100","0000111110001111100011111000","0000101000101010001010100010","0000110101011101010111010101","0000110010111100101111001011","0000111100101111001011110010","0000110111111101111111011111","0000101100011011000110110001","0000011110110111101101111011","0000010010010100100101001001","0000010110000101100001011000","0000010111000101110001011100","0000010100000101000001010000","0000001010000010100000101000","0000001010010010100100101001","0000000110100001101000011010","0000000001010000010100000101","0001000000000000000000000000","0000000100010001000100010001","0000001101100011011000110110","0000010100100101001001010010","0000010111010101110101011101","0000001101110011011100110111","0000010110100101101001011010","0000010101100101011001010110","0000010010110100101101001011","0000101001101010011010100110","0000100100001001000010010000","0000101111001011110010111100","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000101110101011101010111010","0000011100100111001001110010","0000011001100110011001100110","0000011001110110011101100111","0000010011000100110001001100","0001000000000000000000000000","0000001000000010000000100000","0000011111110111111101111111","0000101100001011000010110000","0000011111010111110101111101","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000101100111011001110110011","0000111011011110110111101101","0000011011000110110001101100","0000100111111001111110011111","0000001101000011010000110100","0000101100101011001010110010","0000110000111100001111000011","0000110011111100111111001111","0000111010011110100111101001","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111100011111000111110001","0000111111101111111011111110","0000111111011111110111111101","0000111110011111100111111001","0000111101101111011011110110","0000110011011100110111001101","0000100011011000110110001101","0000001101110011011100110111","0000011110110111101101111011","0000100110101001101010011010","0000101101001011010010110100","0000110010101100101011001010","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000110111011101110111011101","0000110110011101100111011001","0000111111001111110011111100","0000111111011111110111111101","0000111010111110101111101011","0000110011011100110111001101","0000111010101110101011101010","0000111101011111010111110101","0000111011001110110011101100","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111100101111001011110010","0000101100111011001110110011","0000011101010111010101110101","0000101011011010110110101101","0000000000110000001100000011","0000110010101100101011001010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000110101011101010111010101","0000100111011001110110011101","0000101001001010010010100100","0000010011100100111001001110","0000100001011000010110000101","0000011010100110101001101010","0000111101111111011111110111","0000110001001100010011000100","0000001010000010100000101000","0000010000010100000101000001","0000011111100111111001111110","0000011101100111011001110110","0000111111011111110111111101","0000101011011010110110101101","0000100000001000000010000000","0000000011100000111000001110","0000100011111000111110001111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111101011111010111110101","0000111100101111001011110010","0000111111111111111111111111","0000101100101011001010110010","0000000000110000001100000011","0000110110101101101011011010","0000101110111011101110111011","0000110110111101101111011011","0000111111011111110111111101","0000111111111111111111111111","0000111011101110111011101110","0000111110011111100111111001","0000111110001111100011111000","0000100110011001100110011001","0000011100010111000101110001","0000010100000101000001010000","0000100111011001110110011101","0000010101010101010101010101","0000011011110110111101101111","0000101010101010101010101010","0000111101001111010011110100","0000100011001000110010001100","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111100011111000111110001","0000111101001111010011110100","0000101011011010110110101101","0000111110001111100011111000","0000111111111111111111111111","0000111011101110111011101110","0000111110101111101011111010","0000111111111111111111111111","0000110111011101110111011101","0000100000111000001110000011","0000110000011100000111000001","0000110101001101010011010100","0000111011011110110111101101","0000110101001101010011010100","0000111111001111110011111100","0000111110001111100011111000","0000111111101111111011111110","0000111100101111001011110010","0000001011100010111000101110","0000011110110111101101111011","0000100111111001111110011111","0000110111001101110011011100","0000100001111000011110000111","0000011111100111111001111110","0000011010110110101101101011","0000001111000011110000111100","0000011111110111111101111111","0000101001111010011110100111","0000110110101101101011011010","0000101011101010111010101110","0000011100010111000101110001","0000001110010011100100111001","0000000010000000100000001000","0000000100010001000100010001","0001000000000000000000000000","0001000000000000000000000000","0000000001100000011000000110","0000001110000011100000111000","0000100010001000100010001000","0000100101111001011110010111","0000100101111001011110010111","0000011111110111111101111111","0000011001100110011001100110","0000010110000101100001011000","0000010010000100100001001000","0000001110000011100000111000","0000001001000010010000100100","0000000011110000111100001111","0000000101000001010000010100","0000000010110000101100001011","0000001101100011011000110110","0000010111110101111101011111","0000101001011010010110100101","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000110011111100111111001111","0000011001100110011001100110","0000010010100100101001001010","0000011111010111110101111101","0000010000110100001101000011","0000000101000001010000010100","0000000001000000010000000100","0000011101110111011101110111","0000101000101010001010100010","0000101101011011010110110101","0000111110101111101011111010","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111110001111100011111000","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000101100111011001110110011","0000110111011101110111011101","0000100110001001100010011000","0000100011111000111110001111","0000010010000100100001001000","0000101001011010010110100101","0000101110101011101010111010","0000101001101010011010100110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000110011101100111011001110","0000000001110000011100000111","0000001100110011001100110011","0000011101100111011001110110","0000010011010100110101001101","0000110000111100001111000011","0000110110111101101111011011","0000111011111110111111101111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101111111011111110111","0000111100001111000011110000","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111000111110001111100011","0000111011101110111011101110","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000110111001101110011011100","0000010111100101111001011110","0000110111001101110011011100","0000001010010010100100101001","0000101000011010000110100001","0000111111101111111011111110","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111011001110110011101100","0000110100011101000111010001","0000110011101100111011001110","0000011111100111111001111110","0000100110011001100110011001","0000011001100110011001100110","0000111000001110000011100000","0000111011001110110011101100","0000011111010111110101111101","0000010001000100010001000100","0000011011010110110101101101","0000101001001010010010100100","0000110110001101100011011000","0000110001111100011111000111","0000100110111001101110011011","0000001100110011001100110011","0000010011000100110001001100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111110001111100011111000","0000111110111111101111111011","0000111110101111101011111010","0000111101101111011011110110","0000000111110001111100011111","0000011110010111100101111001","0000111100011111000111110001","0000100101101001011010010110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000100100011001000110010001","0000011000010110000101100001","0000100010101000101010001010","0000001010010010100100101001","0000011101000111010001110100","0000111000001110000011100000","0000111000001110000011100000","0000100010011000100110001001","0000111010001110100011101000","0000111000101110001011100010","0000111101001111010011110100","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111011101110111011101110","0000111101111111011111110111","0000111110101111101011111010","0000111101111111011111110111","0000111000001110000011100000","0000101101001011010010110100","0000111101001111010011110100","0000101110101011101010111010","0000111110111111101111111011","0000111111111111111111111111","0000101011001010110010101100","0000110000111100001111000011","0000111000001110000011100000","0000111111101111111011111110","0000100101011001010110010101","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000000100000001000000010000","0000100011001000110010001100","0000100111001001110010011100","0000111001101110011011100110","0000110101101101011011010110","0000010000010100000101000001","0000001101100011011000110110","0000001110010011100100111001","0001000000000000000000000000","0000000011100000111000001110","0001000000000000000000000000","0000000000100000001000000010","0000010011110100111101001111","0000000110010001100100011001","0000000010110000101100001011","0000011010100110101001101010","0000101110101011101010111010","0000111011001110110011101100","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111100011111000111110001","0000111001111110011111100111","0000101111111011111110111111","0000100100101001001010010010","0000100001001000010010000100","0000100101101001011010010110","0000001111100011111000111110","0000010100000101000001010000","0000011000110110001101100011","0000001110110011101100111011","0000001110110011101100111011","0000100110011001100110011001","0000111010111110101111101011","0000111111011111110111111101","0000111110111111101111111011","0000111111001111110011111100","0000111001001110010011100100","0000100000001000000010000000","0000010101010101010101010101","0000101000001010000010100000","0000001001000010010000100100","0000001011000010110000101100","0000000100000001000000010000","0000011000000110000001100000","0000100100001001000010010000","0000110111101101111011011110","0000111111101111111011111110","0000111101001111010011110100","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111101111111011111110111","0000111100111111001111110011","0000111110111111101111111011","0000111010111110101111101011","0000101010001010100010101000","0000101100001011000010110000","0000100011111000111110001111","0000100011011000110110001101","0001000000000000000000000000","0000100000001000000010000000","0000101010001010100010101000","0000111100011111000111110001","0000111100001111000011110000","0000111110011111100111111001","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111011001110110011101100","0000111111111111111111111111","0000111100001111000011110000","0000010110010101100101011001","0001000000000000000000000000","0000011010100110101001101010","0000010100110101001101010011","0000011010010110100101101001","0000011001010110010101100101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111001101110011011100110","0000111111001111110011111100","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000111011011110110111101101","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110100101101001011010010","0000101100101011001010110010","0000101000101010001010100010","0000100001001000010010000100","0000010000010100000101000001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000110110011101100111011001","0000110101011101010111010101","0000101101001011010010110100","0000110010111100101111001011","0000100110101001101010011010","0000111101101111011011110110","0000110110011101100111011001","0000100110001001100010011000","0000001101010011010100110101","0000010110000101100001011000","0000110011101100111011001110","0000111001011110010111100101","0000110110101101101011011010","0000101110011011100110111001","0000010011000100110001001100","0000000011000000110000001100","0000111010101110101011101010","0000111101101111011011110110","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0001000000000000000000000000","0000110000111100001111000011","0000111001101110011011100110","0000100011101000111010001110","0000111111111111111111111111","0000111110101111101011111010","0000111011101110111011101110","0000111110101111101011111010","0000111011001110110011101100","0000111111111111111111111111","0000111001101110011011100110","0000111111101111111011111110","0000010110110101101101011011","0000100001001000010010000100","0000001001010010010100100101","0000100001111000011110000111","0000110111101101111011011110","0000101011001010110010101100","0000110100101101001011010010","0000101011011010110110101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111100001111000011110000","0000111111011111110111111101","0000111001111110011111100111","0000111011001110110011101100","0000101111111011111110111111","0000111111111111111111111111","0000110011111100111111001111","0000110011111100111111001111","0000111001001110010011100100","0000110100101101001011010010","0000110100101101001011010010","0000111100001111000011110000","0000110010111100101111001011","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000000010110000101100001011","0000100101111001011110010111","0000100110111001101110011011","0000101001111010011110100111","0000011000100110001001100010","0000001101010011010100110101","0000000011100000111000001110","0000001001110010011100100111","0000001000100010001000100010","0000000110000001100000011000","0000010000100100001001000010","0000011001000110010001100100","0000100011001000110010001100","0000110000001100000011000000","0000111110111111101111111011","0000111110101111101011111010","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111100101111001011110010","0000111111111111111111111111","0000111010011110100111101001","0000101100101011001010110010","0000110011011100110111001101","0000010111000101110001011100","0000010011100100111001001110","0000010011000100110001001100","0000001110110011101100111011","0000011110000111100001111000","0000110010001100100011001000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100001111000011110000","0000101001011010010110100101","0000010111100101111001011110","0000011111100111111001111110","0000001111000011110000111100","0000000101010001010100010101","0000000011110000111100001111","0000001111110011111100111111","0000101010111010101110101011","0000111000101110001011100010","0000111111001111110011111100","0000111100011111000111110001","0000111110001111100011111000","0000111110101111101011111010","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111100001111000011110000","0000111100101111001011110010","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000110000001100000011000000","0000101001111010011110100111","0000011011100110111001101110","0000011111000111110001111100","0000011011000110110001101100","0001000000000000000000000000","0000001001010010010100100101","0000110010111100101111001011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111101011111010111110101","0000111111001111110011111100","0000111110101111101011111010","0000101000001010000010100000","0001000000000000000000000000","0001000000000000000000000000","0000100001011000010110000101","0000100001111000011110000111","0000010001110100011101000111","0000011011100110111001101110","0000110011011100110111001101","0000111100101111001011110010","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111001111110011111100","0000110100011101000111010001","0000110001001100010011000100","0000100010001000100010001000","0000110100011101000111010001","0000000010100000101000001010","0000111000011110000111100001","0000111001101110011011100110","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000111100001111000011110000","0000111000101110001011100010","0000101110011011100110111001","0000110000101100001011000010","0000110000011100000111000001","0000110111001101110011011100","0000101010011010100110101001","0000111010111110101111101011","0000110101101101011011010110","0000100100001001000010010000","0000010111010101110101011101","0000011110100111101001111010","0000110100111101001111010011","0000111111101111111011111110","0000110100001101000011010000","0000110101101101011011010110","0000011010100110101001101010","0000000100110001001100010011","0000110001011100010111000101","0000111101101111011011110110","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110111111101111111011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000100001011000010110000101","0000001010010010100100101001","0000101011001010110010101100","0000110000101100001011000010","0000101011101010111010101110","0000111011001110110011101100","0000111111111111111111111111","0000111100111111001111110011","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111101011111010111110101","0000100111101001111010011110","0000100110001001100010011000","0001000000000000000000000000","0000101000101010001010100010","0000101101001011010010110100","0000101000111010001110100011","0000111101001111010011110100","0000100001101000011010000110","0000111001111110011111100111","0000111110111111101111111011","0000111111111111111111111111","0000111011101110111011101110","0000111100101111001011110010","0000111111111111111111111111","0000110110111101101111011011","0000111001011110010111100101","0000111111111111111111111111","0000111010111110101111101011","0000110110111101101111011011","0000110011001100110011001100","0000011111110111111101111111","0000111000011110000111100001","0000110110101101101011011010","0000101111001011110010111100","0000110100111101001111010011","0000101000101010001010100010","0000111111111111111111111111","0000110110111101101111011011","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111100001111000011110000","0001000000000000000000000000","0000100000111000001110000011","0000101111001011110010111100","0000100111111001111110011111","0000100010111000101110001011","0000010001000100010001000100","0000010011100100111001001110","0000010100100101001001010010","0000001111110011111100111111","0000010011110100111101001111","0000101010001010100010101000","0000111011011110110111101101","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111111101111111011111110","0000111100001111000011110000","0000111100111111001111110011","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111000001110000011100000","0000110000001100000011000000","0000011111000111110001111100","0000011100010111000101110001","0000010011010100110101001101","0000101001111010011110100111","0000100101111001011110010111","0000110101011101010111010101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000110100011101000111010001","0000100001011000010110000101","0000011100100111001001110010","0000011101010111010101110101","0000001001100010011000100110","0001000000000000000000000000","0000001110110011101100111011","0000100001011000010110000101","0000111011101110111011101110","0000111001101110011011100110","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111101101111011011110110","0000111101001111010011110100","0000111100011111000111110001","0000111100001111000011110000","0000111111101111111011111110","0000111100111111001111110011","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000110010001100100011001000","0000100101111001011110010111","0000011010000110100001101000","0000001101110011011100110111","0000100110001001100010011000","0000001101100011011000110110","0000001101010011010100110101","0000100100001001000010010000","0000110001111100011111000111","0000111010101110101011101010","0000111111111111111111111111","0000111101011111010111110101","0000111100101111001011110010","0000111101101111011011110110","0000101110011011100110111001","0000010111000101110001011100","0000000100010001000100010001","0000010001110100011101000111","0000100001111000011110000111","0000101011001010110010101100","0000011010000110100001101000","0000010010110100101101001011","0000010110000101100001011000","0000011110010111100101111001","0000011011010110110101101101","0000100110011001100110011001","0000100111111001111110011111","0000101101001011010010110100","0000110001101100011011000110","0000111000101110001011100010","0000111010111110101111101011","0000111110011111100111111001","0000111111001111110011111100","0000111000111110001111100011","0000111100111111001111110011","0000111111111111111111111111","0000111100011111000111110001","0000111110101111101011111010","0000111100011111000111110001","0000101101111011011110110111","0000101100011011000110110001","0000100000101000001010000010","0000010110010101100101011001","0000011001010110010101100101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000110100011101000111010001","0000110101101101011011010110","0000111001111110011111100111","0000111100011111000111110001","0000110011011100110111001101","0000111110111111101111111011","0000111011101110111011101110","0000100010011000100110001001","0000100100001001000010010000","0000100111111001111110011111","0000111000011110000111100001","0000111110101111101011111010","0000101101011011010110110101","0000110101111101011111010111","0000011011010110110101101101","0000010000110100001101000011","0000100010101000101010001010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000010100110101001101010011","0000010101000101010001010100","0000101101011011010110110101","0000101100001011000010110000","0000101111001011110010111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000101101011011010110110101","0000110000101100001011000010","0000001011110010111100101111","0000100011111000111110001111","0000101011101010111010101110","0000011111100111111001111110","0000101000011010000110100001","0000110100101101001011010010","0000100011101000111010001110","0000110010101100101011001010","0000111100111111001111110011","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111100101111001011110010","0000110010111100101111001011","0000110110101101101011011010","0000111111111111111111111111","0000101111101011111010111110","0000101110111011101110111011","0000101111111011111110111111","0000101011101010111010101110","0000111001011110010111100101","0000111000001110000011100000","0000100101101001011010010110","0000101010111010101110101011","0000111011001110110011101100","0000110110011101100111011001","0000111111001111110011111100","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0001000000000000000000000000","0000011100000111000001110000","0000110110011101100111011001","0000101011101010111010101110","0000011010000110100001101000","0000100010101000101010001010","0000011111110111111101111111","0000100001111000011110000111","0000100110001001100010011000","0000110100001101000011010000","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000101110011011100110111001","0000100001001000010010000100","0000011011010110110101101101","0000011110000111100001111000","0000100111111001111110011111","0000101111101011111010111110","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111010001110100011101000","0000101100001011000010110000","0000100011011000110110001101","0000011011010110110101101101","0000001110100011101000111010","0000001010000010100000101000","0000001110100011101000111010","0000011110000111100001111000","0000111001101110011011100110","0000111000011110000111100001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111110011111100111111001","0000111111011111110111111101","0000111110111111101111111011","0000111110001111100011111000","0000111101001111010011110100","0000111100001111000011110000","0000111011001110110011101100","0000111010011110100111101001","0000111001111110011111100111","0000111111111111111111111111","0000110001001100010011000100","0000111110111111101111111011","0000111101101111011011110110","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111000011110000111100001","0000101010111010101110101011","0000011100000111000001110000","0000011011100110111001101110","0000011011010110110101101101","0000011010110110101101101011","0000000010110000101100001011","0000010010010100100101001001","0000101011111010111110101111","0000100110101001101010011010","0000110101001101010011010100","0000111100001111000011110000","0000110110101101101011011010","0000100100101001001010010010","0000010110100101101001011010","0000010010010100100101001001","0000001010000010100000101000","0000100000001000000010000000","0000100010101000101010001010","0000011110000111100001111000","0000010000100100001001000010","0000010100110101001101010011","0000010101000101010001010100","0000010100010101000101010001","0000100000101000001010000010","0000011100110111001101110011","0000011101010111010101110101","0000100110001001100010011000","0000101100001011000010110000","0000111000101110001011100010","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000110001001100010011000100","0000111000101110001011100010","0000111101011111010111110101","0000111111001111110011111100","0000111110101111101011111010","0000101101011011010110110101","0000100011011000110110001101","0000100001101000011010000110","0001000000000000000000000000","0000110010101100101011001010","0000111101001111010011110100","0000111100001111000011110000","0000111111111111111111111111","0000111100101111001011110010","0000111111001111110011111100","0000111111101111111011111110","0000111111001111110011111100","0000110011001100110011001100","0000101110001011100010111000","0000111000011110000111100001","0000110101111101011111010111","0000110110111101101111011011","0000111111111111111111111111","0000111111101111111011111110","0000011111010111110101111101","0000100010011000100110001001","0000100101011001010110010101","0000111111111111111111111111","0000111011101110111011101110","0000101001101010011010100110","0000110000001100000011000000","0000010001100100011001000110","0000010101100101011001010110","0000010001110100011101000111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000000100100001001000010010","0000011111010111110101111101","0000100101101001011010010110","0000101011111010111110101111","0000110101011101010111010101","0000111111111111111111111111","0000111110101111101011111010","0000111100101111001011110010","0000111111111111111111111111","0000111011001110110011101100","0000111110011111100111111001","0000111100001111000011110000","0000111111011111110111111101","0000110100111101001111010011","0000110101101101011011010110","0000001110010011100100111001","0000010101010101010101010101","0000110011101100111011001110","0000010111010101110101011101","0000100000011000000110000001","0000101000101010001010100010","0000101100001011000010110000","0000100110101001101010011010","0000100000111000001110000011","0000110010101100101011001010","0000111100101111001011110010","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000110101011101010111010101","0000110010001100100011001000","0000111011001110110011101100","0000101010001010100010101000","0000101100011011000110110001","0000110100001101000011010000","0000110001111100011111000111","0000110000011100000111000001","0000110001101100011011000110","0000100010101000101010001010","0000101010011010100110101001","0000111010101110101011101010","0000111111101111111011111110","0000111111111111111111111111","0000111011011110110111101101","0000111100101111001011110010","0000001001000010010000100100","0000011100010111000101110001","0000101011001010110010101100","0000100111011001110110011101","0000101010101010101010101010","0000101011101010111010101110","0000101110111011101110111011","0000011110110111101101111011","0000110011011100110111001101","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000101011101010111010101110","0000011100110111001101110011","0000011011010110110101101101","0000101000101010001010100010","0000110110111101101111011011","0000111101111111011111110111","0000111111111111111111111111","0000111100001111000011110000","0000111101011111010111110101","0000111100001111000011110000","0000100001101000011010000110","0000011011010110110101101101","0000010101010101010101010101","0000001010010010100100101001","0000000100010001000100010001","0000011111110111111101111111","0000100100001001000010010000","0000110000111100001111000011","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111110011111100111111001","0000111110011111100111111001","0000111101001111010011110100","0000111010101110101011101010","0000110111011101110111011101","0000111110011111100111111001","0000110101001101010011010100","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000101100111011001110110011","0000110110001101100011011000","0000110001001100010011000100","0000111100001111000011110000","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000111101111111011111110111","0000111010101110101011101010","0000100000011000000110000001","0000011100010111000101110001","0000010101010101010101010101","0000101100101011001010110010","0000100001111000011110000111","0000000101000001010000010100","0000000010010000100100001001","0000101011111010111110101111","0000110011001100110011001100","0000100100101001001010010010","0000101010011010100110101001","0000010000010100000101000001","0000011010100110101001101010","0000001010010010100100101001","0000001011100010111000101110","0000100110111001101110011011","0000011111010111110101111101","0000011101000111010001110100","0000010011110100111101001111","0000010010010100100101001001","0000010110000101100001011000","0000001111010011110100111101","0000000101100001011000010110","0000010001100100011001000110","0000001100100011001000110010","0000001011000010110000101100","0000010000010100000101000001","0000010110110101101101011011","0000011110010111100101111001","0000101001001010010010100100","0000110011001100110011001100","0000111100111111001111110011","0000111101011111010111110101","0000101111001011110010111100","0000101011111010111110101111","0000111111111111111111111111","0000111110111111101111111011","0000110111101101111011011110","0000011100010111000101110001","0000010010000100100001001000","0000011110010111100101111001","0000101100111011001110110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110100011101000111010001","0000111111101111111011111110","0000111101011111010111110101","0000111010001110100011101000","0000101000011010000110100001","0000110011101100111011001110","0000111110011111100111111001","0000111010111110101111101011","0000111111111111111111111111","0000111111101111111011111110","0000100101011001010110010101","0000100100001001000010010000","0000101101011011010110110101","0000111111101111111011111110","0000110110111101101111011011","0000100111101001111010011110","0000100001111000011110000111","0000001111100011111000111110","0000011010010110100101101001","0000000000100000001000000010","0000111101101111011011110110","0000111110011111100111111001","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000110110001101100011011000","0000000001110000011100000111","0000100001001000010010000100","0000101000011010000110100001","0000101111001011110010111100","0000101110001011100010111000","0000111011101110111011101110","0000111111101111111011111110","0000111101011111010111110101","0000111111011111110111111101","0000111101001111010011110100","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000110111011101110111011101","0000110111011101110111011101","0000011100010111000101110001","0000001001000010010000100100","0000110001001100010011000100","0000100111001001110010011100","0000010010010100100101001001","0000011010010110100101101001","0000100000011000000110000001","0000100100011001000110010001","0000101001111010011110100111","0000011110010111100101111001","0000100111001001110010011100","0000101001111010011110100111","0000101111001011110010111100","0000101111001011110010111100","0000101010101010101010101010","0000100111101001111010011110","0000101101001011010010110100","0000111001011110010111100101","0000100110101001101010011010","0000100000101000001010000010","0000011011100110111001101110","0000100001111000011110000111","0000100110101001101010011010","0000101111111011111110111111","0000100110011001100110011001","0000101011001010110010101100","0000111010101110101011101010","0000111111111111111111111111","0000110001001100010011000100","0000111100001111000011110000","0000010110110101101101011011","0000010100010101000101010001","0000011110100111101001111010","0000110111111101111111011111","0000101110101011101010111010","0000110010011100100111001001","0000101001001010010010100100","0000101000001010000010100000","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111110111111101111111011","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111110011111100111111001","0000110110011101100111011001","0000101000111010001110100011","0000100000101000001010000010","0000101010011010100110101001","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111110101111101011111010","0000100111101001111010011110","0000011111100111111001111110","0000001101010011010100110101","0000010010110100101101001011","0001000000000000000000000000","0000100011011000110110001101","0000100100111001001110010011","0000101100001011000010110000","0000111111111111111111111111","0000111101111111011111110111","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011111110111111101111","0000111110011111100111111001","0000111100101111001011110010","0000110100001101000011010000","0000110111011101110111011101","0000111000111110001111100011","0000111111111111111111111111","0000111001101110011011100110","0000110111001101110011011100","0000101111001011110010111100","0000111010001110100011101000","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111100101111001011110010","0000111101111111011111110111","0000110001001100010011000100","0000001111110011111100111111","0000100011111000111110001111","0000011111010111110101111101","0000101001101010011010100110","0000010010110100101101001011","0001000000000000000000000000","0000011110000111100001111000","0000110100111101001111010011","0000011001010110010101100101","0000010110010101100101011001","0000010011010100110101001101","0000010101010101010101010101","0000010110000101100001011000","0000100111101001111010011110","0000011000000110000001100000","0000010010100100101001001010","0001000000000000000000000000","0000000001100000011000000110","0000001110010011100100111001","0000010110110101101101011011","0000000101000001010000010100","0000000101100001011000010110","0000010000110100001101000011","0000010111100101111001011110","0000010101010101010101010101","0000010100110101001101010011","0000010110010101100101011001","0000001111000011110000111100","0000000011000000110000001100","0000001011000010110000101100","0000011101010111010101110101","0000101010111010101110101011","0000111010011110100111101001","0000100011101000111010001110","0000110011101100111011001110","0000111000101110001011100010","0000101000011010000110100001","0000001010000010100000101000","0000011011100110111001101110","0000101100111011001110110011","0000111110111111101111111011","0000111101101111011011110110","0000111111011111110111111101","0000111100001111000011110000","0000110010101100101011001010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000100100011001000110010001","0000110011001100110011001100","0000110000011100000111000001","0000111101001111010011110100","0000111111011111110111111101","0000111100001111000011110000","0000110010111100101111001011","0000100001101000011010000110","0000111111111111111111111111","0000111111111111111111111111","0000101011001010110010101100","0000100001011000010110000101","0000011010110110101101101011","0000100000101000001010000010","0000010010100100101001001010","0000000011100000111000001110","0000110100001101000011010000","0000111101011111010111110101","0000111101111111011111110111","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000101101101011011010110110","0001000000000000000000000000","0000011001110110011101100111","0000101001001010010010100100","0000110000111100001111000011","0000100010111000101110001011","0000111011101110111011101110","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000110110101101101011011010","0000111010001110100011101000","0000111110111111101111111011","0000111111111111111111111111","0000110111001101110011011100","0000111011001110110011101100","0000101100011011000110110001","0000100110111001101110011011","0000000001010000010100000101","0000111010101110101011101010","0000101101001011010010110100","0000010111000101110001011100","0000010000110100001101000011","0000010010000100100001001000","0000011101000111010001110100","0000100100011001000110010001","0000010011110100111101001111","0000011001010110010101100101","0000011101100111011001110110","0000011011000110110001101100","0000011011010110110101101101","0000011001110110011101100111","0000010100010101000101010001","0000010110100101101001011010","0000101001101010011010100110","0000011111110111111101111111","0000100100011001000110010001","0000100111111001111110011111","0000100111111001111110011111","0000100100011001000110010001","0000100001111000011110000111","0000100101001001010010010100","0000100101101001011010010110","0000111010011110100111101001","0000101101101011011010110110","0000101101001011010010110100","0000011000110110001101100011","0000000110000001100000011000","0000100001101000011010000110","0000110000101100001011000010","0000111101001111010011110100","0000110000001100000011000000","0000101001111010011110100111","0000110100101101001011010010","0000111111101111111011111110","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111111111111111111111111","0000111101011111010111110101","0000111100101111001011110010","0000111111111111111111111111","0000111111001111110011111100","0000110011111100111111001111","0000101000011010000110100001","0000101011111010111110101111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101110011011100110111001","0000110011101100111011001110","0000000000110000001100000011","0000011110110111101101111011","0000000010110000101100001011","0000010111110101111101011111","0000011111100111111001111110","0000011011010110110101101101","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111001101110011011100110","0000111100111111001111110011","0000111101001111010011110100","0000111001101110011011100110","0000110000111100001111000011","0000111111111111111111111111","0000111001011110010111100101","0000101100001011000010110000","0000110001101100011011000110","0000110110111101101111011011","0000110011011100110111001101","0000110011111100111111001111","0000100101101001011010010110","0000111001001110010011100100","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000110101001101010011010100","0000100001111000011110000111","0000100101101001011010010110","0000011000010110000101100001","0000101001111010011110100111","0000011111000111110001111100","0000000000110000001100000011","0000011111000111110001111100","0000100000011000000110000001","0000100011111000111110001111","0000010010000100100001001000","0000010101110101011101010111","0000011011000110110001101100","0000000101010001010100010101","0001000000000000000000000000","0000001110000011100000111000","0000010110000101100001011000","0000010011000100110001001100","0000011010010110100101101001","0000101001001010010010100100","0000101101101011011010110110","0000110011111100111111001111","0000101011011010110110101101","0000100101011001010110010101","0000100100011001000110010001","0000100001111000011110000111","0000011110000111100001111000","0000100000011000000110000001","0000100110111001101110011011","0000010101110101011101010111","0000001001010010010100100101","0000000010110000101100001011","0000000111010001110100011101","0000100110011001100110011001","0000101010101010101010101010","0000100111111001111110011111","0000011110110111101101111011","0000001000100010001000100010","0000001111010011110100111101","0000100011111000111110001111","0000111111111111111111111111","0000111110111111101111111011","0000110010001100100011001000","0000110001011100010111000101","0000111001011110010111100101","0000111011001110110011101100","0000111111001111110011111100","0000111111111111111111111111","0000100101011001010110010101","0000110101111101011111010111","0000100110011001100110011001","0000111111111111111111111111","0000111110011111100111111001","0000111101011111010111110101","0000111010001110100011101000","0000101100111011001110110011","0000111111111111111111111111","0000111110001111100011111000","0000101011101010111010101110","0000011100000111000001110000","0000001101100011011000110110","0000100011101000111010001110","0000000111100001111000011110","0000010001100100011001000110","0000100110011001100110011001","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000101111001011110010111100","0000000000010000000100000001","0000010011000100110001001100","0000011011010110110101101101","0000011110000111100001111000","0000101100011011000110110001","0000110001101100011011000110","0000111110111111101111111011","0000111111101111111011111110","0000111110011111100111111001","0000101111011011110110111101","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111101011111010111110101","0000100000001000000010000000","0000110110111101101111011011","0000100101101001011010010110","0001000000000000000000000000","0000101000011010000110100001","0000110100111101001111010011","0000101011101010111010101110","0000011110010111100101111001","0000011110100111101001111010","0000011011010110110101101101","0000011101000111010001110100","0000011110000111100001111000","0000100011101000111010001110","0000101101001011010010110100","0000100010011000100110001001","0000010110000101100001011000","0000011110100111101001111010","0000100001101000011010000110","0000110011011100110111001101","0000101011011010110110101101","0000100100101001001010010010","0000101001011010010110100101","0000101110011011100110111001","0000100001001000010010000100","0000100001111000011110000111","0000010101100101011001010110","0000011110100111101001111010","0000011011110110111101101111","0000011100100111001001110010","0000100100111001001110010011","0000101010111010101110101011","0000000010000000100000001000","0000101011001010110010101100","0000100111111001111110011111","0000111001101110011011100110","0000101111011011110110111101","0000101100101011001010110010","0000111000101110001011100010","0000111101101111011011110110","0000111100101111001011110010","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111010111110101111101011","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000101111111011111110111111","0000101101001011010010110100","0000111111001111110011111100","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000101111011011110110111101","0001000000000000000000000000","0000010110100101101001011010","0000010010010100100101001001","0000001001010010010100100101","0000010001110100011101000111","0000011111010111110101111101","0000110001101100011011000110","0000110011011100110111001101","0000111000011110000111100001","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111001001110010011100100","0000110011111100111111001111","0000110001001100010011000100","0000110100101101001011010010","0000011100010111000101110001","0000100010001000100010001000","0000100100011001000110010001","0000100011111000111110001111","0000010110000101100001011000","0000101011101010111010101110","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111110111111101111111011","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111011001110110011101100","0000101110001011100010111000","0000111010011110100111101001","0000100110001001100010011000","0000100110001001100010011000","0000101100111011001110110011","0000000010100000101000001010","0000100011011000110110001101","0000100100011001000110010001","0000010000110100001101000011","0001000000000000000000000000","0000010011000100110001001100","0000010011110100111101001111","0000001100110011001100110011","0000010000100100001001000010","0000011100000111000001110000","0000011000100110001001100010","0000100011011000110110001101","0000110010001100100011001000","0000111111001111110011111100","0000111111111111111111111111","0000111101001111010011110100","0000111001101110011011100110","0000110101101101011011010110","0000110000001100000011000000","0000101010001010100010101000","0000100101111001011110010111","0000100100101001001010010010","0000100001101000011010000110","0000100000111000001110000011","0000101100011011000110110001","0000011011100110111001101110","0000000010100000101000001010","0000000101110001011100010111","0000010111100101111001011110","0000011010010110100101101001","0000000010010000100100001001","0000001100100011001000110010","0000011010110110101101101011","0000100101111001011110010111","0000100101111001011110010111","0000100110011001100110011001","0000101101111011011110110111","0000110110001101100011011000","0000110010001100100011001000","0000111010101110101011101010","0000111111111111111111111111","0000101110011011100110111001","0000111010011110100111101001","0000101011101010111010101110","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000110101101101011011010110","0000111011001110110011101100","0000111111111111111111111111","0000111101101111011011110110","0000010111000101110001011100","0000010010110100101101001011","0000010100100101001001010010","0000100111101001111010011110","0000000101000001010000010100","0000011100010111000101110001","0000010010110100101101001011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000110010111100101111001011","0000000100000001000000010000","0000001001010010010100100101","0000011101000111010001110100","0000100011111000111110001111","0000010010000100100001001000","0000101110111011101110111011","0000111111111111111111111111","0000111010011110100111101001","0000111011001110110011101100","0000101010101010101010101010","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111101011111010111110101","0000111010111110101111101011","0000100001101000011010000110","0000111110011111100111111001","0000111101101111011011110110","0000100100111001001110010011","0001000000000000000000000000","0000001110100011101000111010","0000011010000110100001101000","0000011010110110101101101011","0000010100010101000101010001","0000100101011001010110010101","0000110001011100010111000101","0000110101111101011111010111","0000110111001101110011011100","0000110011101100111011001110","0000101001001010010010100100","0000100110101001101010011010","0000100100101001001010010010","0000010001110100011101000111","0000010100110101001101010011","0000100101011001010110010101","0000011011110110111101101111","0000011011000110110001101100","0000010010010100100101001001","0000010010110100101101001011","0000010111100101111001011110","0000010011000100110001001100","0000001001110010011100100111","0000010101110101011101010111","0000101101001011010010110100","0000101011011010110110101101","0000101010111010101110101011","0000000010000000100000001000","0000011110100111101001111010","0000110100101101001011010010","0000100111111001111110011111","0000110011111100111111001111","0000110010111100101111001011","0000101111111011111110111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000110011101100111011001110","0000111001101110011011100110","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111011101110111011101110","0000110101011101010111010101","0000110000111100001111000011","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110011001100110011001100","0000100001001000010010000100","0001000000000000000000000000","0000010100000101000001010000","0000010110110101101101011011","0000000000010000000100000001","0000001101100011011000110110","0000011011010110110101101101","0000100101111001011110010111","0000111110001111100011111000","0000111001001110010011100100","0000110111001101110011011100","0000111010011110100111101001","0000111100101111001011110010","0000111010111110101111101011","0000111010001110100011101000","0000111011101110111011101110","0000110111101101111011011110","0000101110001011100010111000","0000100000101000001010000010","0000011111010111110101111101","0000010111110101111101011111","0000010110000101100001011000","0000010100100101001001010010","0000011101000111010001110100","0000010111100101111001011110","0000011110010111100101111001","0000111000111110001111100011","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111100011111000111110001","0000111111111111111111111111","0000111010011110100111101001","0000111010111110101111101011","0000111001101110011011100110","0000111000011110000111100001","0000101101001011010010110100","0000101010111010101110101011","0000010001000100010001000100","0000001100010011000100110001","0000001111110011111100111111","0000001001010010010100100101","0000010001100100011001000110","0000011010010110100101101001","0000010010100100101001001010","0000010010010100100101001001","0000011011100110111001101110","0000100101101001011010010110","0000101111011011110110111101","0000101011111010111110101111","0000110101111101011111010111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111001001110010011100100","0000110010011100100111001001","0000101010011010100110101001","0000011111010111110101111101","0000100011011000110110001101","0000011111100111111001111110","0000011000100110001001100010","0000000001000000010000000100","0000000111100001111000011110","0000010100000101000001010000","0000011111110111111101111111","0000100011011000110110001101","0000010110100101101001011010","0000010010000100100001001000","0000011100100111001001110010","0000101101011011010110110101","0000111000011110000111100001","0000110001011100010111000101","0000111001011110010111100101","0000111110001111100011111000","0000111000011110000111100001","0000111010111110101111101011","0000111000101110001011100010","0000111110111111101111111011","0000111111011111110111111101","0000111101111111011111110111","0000111010001110100011101000","0000111101101111011011110110","0000111111111111111111111111","0000110111011101110111011101","0000001001000010010000100100","0000010000010100000101000001","0000010110000101100001011000","0000110010101100101011001010","0000001111010011110100111101","0000011101010111010101110101","0001000000000000000000000000","0000111111001111110011111100","0000111110001111100011111000","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000101010111010101110101011","0000001000000010000000100000","0000101000011010000110100001","0000001111010011110100111101","0000100001111000011110000111","0000100011011000110110001101","0000100011101000111010001110","0000110101101101011011010110","0000110111101101111011011110","0000111100101111001011110010","0000100111101001111010011110","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111111001111110011111100","0000110001101100011011000110","0000100010111000101110001011","0000100000011000000110000001","0000001100100011001000110010","0000000011110000111100001111","0000000011110000111100001111","0001000000000000000000000000","0000000100100001001000010010","0001000000000000000000000000","0001000000000000000000000000","0000000010000000100000001000","0000000010000000100000001000","0000000110000001100000011000","0000011010100110101001101010","0000100011011000110110001101","0000100100101001001010010010","0000100001101000011010000110","0000010010100100101001001010","0000001110100011101000111010","0000001011110010111100101111","0000010010100100101001001010","0000001111000011110000111100","0000001010000010100000101000","0000001010100010101000101010","0000010000100100001001000010","0000010011110100111101001111","0000010101000101010001010100","0000001100110011001100110011","0000001100100011001000110010","0000010111110101111101011111","0000100001011000010110000101","0000101110101011101010111010","0000011000000110000001100000","0000000000010000000100000001","0000101110111011101110111011","0000101010101010101010101010","0000101101101011011010110110","0000111111111111111111111111","0000101000001010000010100000","0000111010111110101111101011","0000111110111111101111111011","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111010011110100111101001","0000101100101011001010110010","0000110001001100010011000100","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111001001110010011100100","0000110110111101101111011011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110001011100010111000101","0000011101000111010001110100","0000001110010011100100111001","0000000110110001101100011011","0000010011100100111001001110","0000000111110001111100011111","0001000000000000000000000000","0000011011010110110101101101","0000100100011001000110010001","0000101110111011101110111011","0000110101001101010011010100","0000111000011110000111100001","0000110101111101011111010111","0000110010101100101011001010","0000110001001100010011000100","0000101101111011011110110111","0000101001101010011010100110","0000101000011010000110100001","0000100000101000001010000010","0000011110000111100001111000","0000001111110011111100111111","0000010010100100101001001010","0000001011110010111100101111","0000010011000100110001001100","0000010001110100011101000111","0000100110101001101010011010","0000011100100111001001110010","0000110010011100100111001001","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111001001110010011100100","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000110011011100110111001101","0000110000001100000011000000","0000101100001011000010110000","0000010100110101001101010011","0000000101000001010000010100","0000001010100010101000101010","0000010011010100110101001101","0000011100010111000101110001","0000000101000001010000010100","0000100010001000100010001000","0000011111010111110101111101","0000011011110110111101101111","0000101010101010101010101010","0000111001001110010011100100","0000111001111110011111100111","0000110111111101111111011111","0000111011111110111111101111","0000111111011111110111111101","0000111101001111010011110100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111111101111111011111110","0000111101101111011011110110","0000111011111110111111101111","0000110011011100110111001101","0000100001001000010010000100","0000101001011010010110100101","0000101000011010000110100001","0000100110111001101110011011","0000101110101011101010111010","0000101010011010100110101001","0000011110000111100001111000","0000011000000110000001100000","0000011000100110001001100010","0000100101011001010110010101","0000101010111010101110101011","0000110000011100000111000001","0000111000101110001011100010","0000111001001110010011100100","0000111100101111001011110010","0000111101011111010111110101","0000111101101111011011110110","0000111001001110010011100100","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111101111111011111110111","0000111111101111111011111110","0000111011001110110011101100","0000101000001010000010100000","0000010011110100111101001111","0000001101000011010000110100","0000010011100100111001001110","0000100111111001111110011111","0000011100100111001001110010","0000100000011000000110000001","0001000000000000000000000000","0000110010011100100111001001","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000010101100101011001010110","0000001010000010100000101000","0000110101001101010011010100","0000011011010110110101101101","0000011111100111111001111110","0000100010101000101010001010","0000101001011010010110100101","0000100011011000110110001101","0000110011111100111111001111","0000110101001101010011010100","0000101100011011000110110001","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111011101110111011101110","0000011011000110110001101100","0000001000100010001000100010","0001000000000000000000000000","0000001110010011100100111001","0000011011000110110001101100","0000101000001010000010100000","0000100011101000111010001110","0000011101110111011101110111","0000011101000111010001110100","0000100010001000100010001000","0000100000011000000110000001","0000010110110101101101011011","0000001010010010100100101001","0000001100010011000100110001","0000000011010000110100001101","0000000001100000011000000110","0000010001010100010101000101","0000010100000101000001010000","0000010100000101000001010000","0000001111100011111000111110","0000001000110010001100100011","0000001011100010111000101110","0000001100110011001100110011","0000010001000100010001000100","0000001010110010101100101011","0000010001110100011101000111","0000010000010100000101000001","0000001101010011010100110101","0000001010110010101100101011","0000001101000011010000110100","0000001101010011010100110101","0000011100110111001101110011","0000100101001001010010010100","0000000100000001000000010000","0000010000100100001001000010","0000101010111010101110101011","0000100111011001110110011101","0000111100101111001011110010","0000110001011100010111000101","0000101111111011111110111111","0000111111011111110111111101","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111110011111100111111001","0000111000001110000011100000","0000100111111001111110011111","0000101110011011100110111001","0000111101011111010111110101","0000111100111111001111110011","0000111110011111100111111001","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000111011011110110111101101","0000111010111110101111101011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000101100011011000110110001","0000100010101000101010001010","0000001111110011111100111111","0000001011010010110100101101","0000001110000011100000111000","0000001100010011000100110001","0000001000110010001100100011","0000010110000101100001011000","0000100111101001111010011110","0000101010101010101010101010","0000110001011100010111000101","0000110000111100001111000011","0000100111111001111110011111","0000100100001001000010010000","0000100110111001101110011011","0000100100101001001010010010","0000011101010111010101110101","0000011101000111010001110100","0000100001001000010010000100","0000011000110110001101100011","0000010110100101101001011010","0000010011000100110001001100","0000001101010011010100110101","0000001001100010011000100110","0000010111110101111101011111","0000101001101010011010100110","0000100011111000111110001111","0000110100101101001011010010","0000111111111111111111111111","0000111100111111001111110011","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000110010001100100011001000","0000010110000101100001011000","0000010010110100101101001011","0000000000010000000100000001","0000001101010011010100110101","0000010000110100001101000011","0000010011010100110101001101","0000011010100110101001101010","0000100010001000100010001000","0000110010011100100111001001","0000101101011011010110110101","0000110001001100010011000100","0000101010111010101110101011","0000111000111110001111100011","0000111011001110110011101100","0000111100111111001111110011","0000111110001111100011111000","0000111110111111101111111011","0000111110111111101111111011","0000111110011111100111111001","0000111110011111100111111001","0000111111011111110111111101","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111010001110100011101000","0000110111101101111011011110","0000111101011111010111110101","0000111000111110001111100011","0000110111001101110011011100","0000111001111110011111100111","0000110011011100110111001101","0000110101111101011111010111","0000110001001100010011000100","0000110001101100011011000110","0000111010011110100111101001","0000111110011111100111111001","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111010101110101011101010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000110010101100101011001010","0000011111100111111001111110","0000010100100101001001010010","0000001110110011101100111011","0000011111110111111101111111","0000011011010110110101101101","0000100010111000101110001011","0000011101100111011001110110","0000010010010100100101001001","0000100011001000110010001100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000000010000000100000001000","0000001010100010101000101010","0000101101101011011010110110","0000101110001011100010111000","0000001100010011000100110001","0000100010111000101110001011","0000101101001011010010110100","0000010101010101010101010101","0000100101101001011010010110","0000101101001011010010110100","0000110100011101000111010001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000100000011000000110000001","0000000000100000001000000010","0000001000000010000000100000","0000110001101100011011000110","0000111100101111001011110010","0000111100101111001011110010","0000110111011101110111011101","0000111010001110100011101000","0000111010101110101011101010","0000111011101110111011101110","0000110111011101110111011101","0000101111101011111010111110","0000101001011010010110100101","0000100000101000001010000010","0000101101011011010110110101","0000101101111011011110110111","0000010001010100010101000101","0000001101110011011100110111","0000100000111000001110000011","0000100001001000010010000100","0000011000100110001001100010","0000011010010110100101101001","0000010110110101101101011011","0000100111101001111010011110","0000011110000111100001111000","0000010110100101101001011010","0000011110110111101101111011","0000010011100100111001001110","0000011011100110111001101110","0000010001110100011101000111","0000011111100111111001111110","0000011000100110001001100010","0000001011110010111100101111","0000000111010001110100011101","0000001011100010111000101110","0001000000000000000000000000","0000010100110101001101010011","0000101101001011010010110100","0000100011111000111110001111","0000111111111111111111111111","0000110111111101111111011111","0000111101011111010111110101","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111110101111101011111010","0000111010111110101111101011","0000111100111111001111110011","0000110111001101110011011100","0000100101111001011110010111","0000110001001100010011000100","0000111011001110110011101100","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111101111111011111110111","0000111100101111001011110010","0000111011111110111111101111","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111100111111001111110011","0000111101011111010111110101","0000111101101111011011110110","0000100111001001110010011100","0000100101101001011010010110","0000011010000110100001101000","0000011001100110011001100110","0000010011100100111001001110","0000001100110011001100110011","0000010101100101011001010110","0000010100110101001101010011","0000010100000101000001010000","0000100011101000111010001110","0000011100010111000101110001","0000011010110110101101101011","0000100100001001000010010000","0000101111001011110010111100","0000110000111100001111000011","0000101010001010100010101000","0000100011101000111010001110","0000011000100110001001100010","0000011001010110010101100101","0000011101010111010101110101","0000010100110101001101010011","0000010011000100110001001100","0000011100010111000101110001","0000101000011010000110100001","0000100010101000101010001010","0000101001101010011010100110","0000100111111001111110011111","0000110000001100000011000000","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111001111110011111100","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111111001111110011111100","0000111010011110100111101001","0000110011101100111011001110","0000101000111010001110100011","0000101100011011000110110001","0000100111011001110110011101","0000001100110011001100110011","0000000100010001000100010001","0000010000110100001101000011","0000010110100101101001011010","0000011100010111000101110001","0000101001101010011010100110","0000110001011100010111000101","0000110111111101111111011111","0000111111011111110111111101","0000111010111110101111101011","0000111000101110001011100010","0000111110011111100111111001","0000111110001111100011111000","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111110001111100011111000","0000111111011111110111111101","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111101101111011011110110","0000111011101110111011101110","0000111111111111111111111111","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000011110110111101101111011","0000011111010111110101111101","0000010110000101100001011000","0000100110001001100010011000","0000011101000111010001110100","0000100101011001010110010101","0000100011011000110110001101","0000010001000100010001000100","0000100011111000111110001111","0000011010000110100001101000","0000111110001111100011111000","0000111100101111001011110010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111100101111001011110010","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111100011111000111110001","0000100010111000101110001011","0000000011100000111000001110","0000010110100101101001011010","0000101010011010100110101001","0000111101001111010011110100","0000110101111101011111010111","0000010110000101100001011000","0000110101011101010111010101","0000010100110101001101010011","0000101101011011010110110101","0000101011101010111010101110","0000101101001011010010110100","0000111100011111000111110001","0000111110011111100111111001","0000101101001011010010110100","0000000111010001110100011101","0000010110010101100101011001","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000110010011100100111001001","0000101000001010000010100000","0000011111100111111001111110","0000011010000110100001101000","0000010111010101110101011101","0000010110100101101001011010","0000011011010110110101101101","0000001111110011111100111111","0000010010000100100001001000","0000011011100110111001101110","0000010000000100000001000000","0000010101110101011101010111","0000010010010100100101001001","0000011101010111010101110101","0000100001001000010010000100","0000101001011010010110100101","0000011000110110001101100011","0000000101110001011100010111","0000001010100010101000101010","0000011000100110001001100010","0000001001010010010100100101","0000001101100011011000110110","0000000001110000011100000111","0000010111100101111001011110","0000101010011010100110101001","0000100111011001110110011101","0000111001101110011011100110","0000111011011110110111101101","0000111111111111111111111111","0000111111101111111011111110","0000111100001111000011110000","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111011101110111011101110","0000111110101111101011111010","0000110010011100100111001001","0000110010101100101011001010","0000101101001011010010110100","0000111111111111111111111111","0000110000111100001111000011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111100011111000111110001","0000100010001000100010001000","0000100111011001110110011101","0000011000010110000101100001","0000001100000011000000110000","0000000011110000111100001111","0000001101010011010100110101","0000011000010110000101100001","0000011101000111010001110100","0000010010100100101001001010","0001000000000000000000000000","0000011001110110011101100111","0000100011101000111010001110","0000100111011001110110011101","0000011110010111100101111001","0000011011010110110101101101","0000011001010110010101100101","0000011000010110000101100001","0000100010111000101110001011","0000011100110111001101110011","0000101000101010001010100010","0000100111101001111010011110","0000100011011000110110001101","0000100001101000011010000110","0000100110011001100110011001","0000101001011010010110100101","0000011111000111110001111100","0000100010011000100110001001","0000010001010100010101000101","0000110101111101011111010111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111011001110110011101100","0000110001111100011111000111","0000110101001101010011010100","0000111111111111111111111111","0000111111111111111111111111","0000011000010110000101100001","0000001001100010011000100110","0000001001010010010100100101","0000011010110110101101101011","0000010011100100111001001110","0000100101111001011110010111","0000101101011011010110110101","0000110100101101001011010010","0000111011111110111111101111","0000111110001111100011111000","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111011001110110011101100","0000111101101111011011110110","0000111110001111100011111000","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111111011111110111111101","0000101111111011111110111111","0000101101111011011110110111","0000100111111001111110011111","0000101011011010110110101101","0000101100111011001110110011","0000110011001100110011001100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111101001111010011110100","0000111111001111110011111100","0000101111101011111010111110","0000100000111000001110000011","0000110000011100000111000001","0000011010010110100101101001","0000000110010001100100011001","0000000110010001100100011001","0000001111110011111100111111","0000001001110010011100100111","0000101010101010101010101010","0000100001101000011010000110","0000000011110000111100001111","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000001000100010001000100010","0000001110010011100100111001","0000010000010100000101000001","0000101010111010101110101011","0000100011101000111010001110","0000110100001101000011010000","0000110111001101110011011100","0000011100010111000101110001","0000100010001000100010001000","0000011101010111010101110101","0000110011011100110111001101","0000110100001101000011010000","0000100001111000011110000111","0000110001011100010111000101","0000100001101000011010000110","0000100100101001001010010010","0000111111001111110011111100","0000111110101111101011111010","0000111111011111110111111101","0000111111001111110011111100","0000111110011111100111111001","0000111101111111011111110111","0000111110011111100111111001","0000111111001111110011111100","0000111111011111110111111101","0000111110111111101111111011","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111000111110001111100011","0000110001001100010011000100","0000101001001010010010100100","0000100100001001000010010000","0000010110100101101001011010","0000100000011000000110000001","0000010011100100111001001110","0000010101000101010001010100","0000110101101101011011010110","0000111010111110101111101011","0000100101011001010110010101","0000111101101111011011110110","0000101011111010111110101111","0000101101001011010010110100","0000011100100111001001110010","0000011100010111000101110001","0000001011010010110100101101","0000001010000010100000101000","0000011000100110001001100010","0000010011010100110101001101","0000100000101000001010000010","0000001011100010111000101110","0000010101000101010001010100","0000100000111000001110000011","0000100110111001101110011011","0000101101001011010010110100","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111101011111010111110101","0000111111101111111011111110","0000111101101111011011110110","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000110110111101101111011011","0000110100001101000011010000","0000100111101001111010011110","0000100100111001001110010011","0000100010001000100010001000","0000110100101101001011010010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000100011111000111110001111","0000100000111000001110000011","0000011000000110000001100000","0000000101010001010100010101","0000010000100100001001000010","0000000011000000110000001100","0000001111100011111000111110","0000001101000011010000110100","0000011110000111100001111000","0000100000011000000110000001","0000010000110100001101000011","0000000000110000001100000011","0000000110110001101100011011","0000001011110010111100101111","0000001001100010011000100110","0000001100000011000000110000","0000010111000101110001011100","0000001100000011000000110000","0000001101010011010100110101","0000010011110100111101001111","0000100000101000001010000010","0000011010010110100101101001","0000010011000100110001001100","0000001101010011010100110101","0000001100110011001100110011","0000010011110100111101001111","0000010110100101101001011010","0000010110100101101001011010","0000101001101010011010100110","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111010011110100111101001","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111010001110100011101000","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000100000001000000010000000","0001000000000000000000000000","0000000011000000110000001100","0000010110100101101001011010","0000001111010011110100111101","0000100011001000110010001100","0000101101101011011010110110","0000110101101101011011010110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111001011110010111100101","0000110011101100111011001110","0000100011001000110010001100","0000100101111001011110010111","0000110101011101010111010101","0000110100111101001111010011","0000101011011010110110101101","0000100111011001110110011101","0000110000101100001011000010","0000100110001001100010011000","0000011100010111000101110001","0000101000111010001110100011","0000110000111100001111000011","0000111100011111000111110001","0000111011001110110011101100","0000111101111111011111110111","0000111111001111110011111100","0000111100001111000011110000","0000111110101111101011111010","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000110100111101001111010011","0000101111011011110110111101","0000101111011011110110111101","0000110101101101011011010110","0000000110000001100000011000","0000110010001100100011001000","0000010011110100111101001111","0000010110000101100001011000","0000001000010010000100100001","0000010010010100100101001001","0000100100101001001010010010","0000000000100000001000000010","0000111001011110010111100101","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111011111110111111101","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000110001101100011011000110","0001000000000000000000000000","0000010010010100100101001001","0000010011000100110001001100","0000100100101001001010010010","0000101100001011000010110000","0000101000011010000110100001","0000011101010111010101110101","0000011101110111011101110111","0000000000110000001100000011","0000011011010110110101101101","0000101001111010011110100111","0000111000111110001111100011","0000111111111111111111111111","0000011101010111010101110101","0000011001110110011101100111","0000111111101111111011111110","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111101111111011111110111","0000111100001111000011110000","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111110111111101111111011","0000111100011111000111110001","0000100011001000110010001100","0000101000111010001110100011","0000011011010110110101101101","0000101001001010010010100100","0000101111011011110110111101","0000110010011100100111001001","0000110100101101001011010010","0000111111111111111111111111","0000110000011100000111000001","0000100110101001101010011010","0000010111110101111101011111","0000100000101000001010000010","0000011000010110000101100001","0000011001010110010101100101","0000101011001010110010101100","0000100100111001001110010011","0000100001101000011010000110","0000010010010100100101001001","0000001100100011001000110010","0000011100100111001001110010","0000101000001010000010100000","0000101110011011100110111001","0000110111011101110111011101","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111011101110111011101110","0000111101011111010111110101","0000111011001110110011101100","0000111111111111111111111111","0000111011001110110011101100","0000110110011101100111011001","0000101110101011101010111010","0000100011111000111110001111","0000001001100010011000100110","0000000010110000101100001011","0000010001110100011101000111","0000100101001001010010010100","0000101010111010101110101011","0000101111001011110010111100","0000111111111111111111111111","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000100110011001100110011001","0000100001101000011010000110","0000010111110101111101011111","0000010011110100111101001111","0000010000110100001101000011","0000001000110010001100100011","0000000110010001100100011001","0000010000010100000101000001","0000010111010101110101011101","0000010010100100101001001010","0000001111110011111100111111","0000001001110010011100100111","0001000000000000000000000000","0000000001110000011100000111","0000000010110000101100001011","0000000000010000000100000001","0001000000000000000000000000","0001000000000000000000000000","0000000001000000010000000100","0001000000000000000000000000","0000001100000011000000110000","0000010000000100000001000000","0000010010110100101101001011","0000011011100110111001101110","0000100100011001000110010001","0000100001001000010010000100","0000100010111000101110001011","0000101001011010010110100101","0000101101111011011110110111","0000110110101101101011011010","0000111101101111011011110110","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110000001100000011000000","0000010101010101010101010101","0001000000000000000000000000","0000001100000011000000110000","0000010100000101000001010000","0000010100010101000101010001","0000010110000101100001011000","0000111011001110110011101100","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111110011111100111111001","0000111111011111110111111101","0000111111101111111011111110","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111001001110010011100100","0000111000011110000111100001","0000110010111100101111001011","0000101111101011111010111110","0000011111110111111101111111","0000001110010011100100111001","0000110011111100111111001111","0000101001001010010010100100","0000010101100101011001010110","0000001010010010100100101001","0000001001000010010000100100","0000010110100101101001011010","0000010001000100010001000100","0000011000100110001001100010","0000100000111000001110000011","0000011011010110110101101101","0000011110110111101101111011","0000011001100110011001100110","0000100111011001110110011101","0000111001001110010011100100","0000111111001111110011111100","0000111111111111111111111111","0000111011101110111011101110","0000111001101110011011100110","0000111110111111101111111011","0000111110011111100111111001","0000111011101110111011101110","0000110110111101101111011011","0000111000001110000011100000","0000110011001100110011001100","0000111000011110000111100001","0000010011000100110001001100","0000111001001110010011100100","0000110011101100111011001110","0000101000111010001110100011","0000001100110011001100110011","0000000100110001001100010011","0000000011000000110000001100","0000010011100100111001001110","0000000010000000100000001000","0000101100111011001110110011","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000011111000111110001111100","0000000000100000001000000010","0000010101110101011101010111","0000011100000111000001110000","0000011011010110110101101101","0000100001101000011010000110","0000010111010101110101011101","0000011110010111100101111001","0000100011001000110010001100","0000000101100001011000010110","0000011000110110001101100011","0000110011011100110111001101","0000111111111111111111111111","0000111010101110101011101010","0000110111011101110111011101","0000110100011101000111010001","0000110001101100011011000110","0000111111101111111011111110","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111101011111010111110101","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111101101111011011110110","0000111101101111011011110110","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000110110101101101011011010","0000101011001010110010101100","0000110011101100111011001110","0000101101001011010010110100","0000110100011101000111010001","0000101100001011000010110000","0000110011011100110111001101","0000101011111010111110101111","0000011111100111111001111110","0000010100010101000101010001","0000011111100111111001111110","0000010001000100010001000100","0000001111110011111100111111","0000001110110011101100111011","0000010011010100110101001101","0000010001100100011001000110","0000001010010010100100101001","0000001011010010110100101101","0000001010010010100100101001","0000001111000011110000111100","0000010100100101001001010010","0000100001001000010010000100","0000110001001100010011000100","0000110100001101000011010000","0000111100101111001011110010","0000111110011111100111111001","0000111010001110100011101000","0000111110011111100111111001","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000101111011011110110111101","0000101111011011110110111101","0000011111000111110001111100","0000001011010010110100101101","0000000111100001111000011110","0000010011100100111001001110","0000000000100000001000000010","0000010011010100110101001101","0000101100101011001010110010","0000111010011110100111101001","0000110100111101001111010011","0000110110111101101111011011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000100111111001111110011111","0000011011100110111001101110","0000011001010110010101100101","0000001010100010101000101010","0000001001000010010000100100","0000010000010100000101000001","0000001110100011101000111010","0000001110110011101100111011","0000001000000010000000100000","0000000001000000010000000100","0000000100100001001000010010","0000001101010011010100110101","0000001011000010110000101100","0000011000110110001101100011","0000100001101000011010000110","0000100101011001010110010101","0000101000011010000110100001","0000100100111001001110010011","0000100100011001000110010001","0000011110010111100101111001","0000011001100110011001100110","0000010110010101100101011001","0000000100100001001000010010","0000000111110001111100011111","0000010101000101010001010100","0000010111010101110101011101","0000101000111010001110100011","0000101100111011001110110011","0000111010001110100011101000","0000101110111011101110111011","0000100111101001111010011110","0000111011111110111111101111","0000111101101111011011110110","0000111110111111101111111011","0000111100011111000111110001","0000111111001111110011111100","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111101101111011011110110","0000110100101101001011010010","0000101000001010000010100000","0000100010101000101010001010","0000010010100100101001001010","0000000011000000110000001100","0000010010110100101101001011","0000001111000011110000111100","0000011011110110111101101111","0000101010111010101110101011","0000111010001110100011101000","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111001111110011111100","0000111111101111111011111110","0000110110101101101011011010","0000011001110110011101100111","0000100010011000100110001001","0000100011001000110010001100","0000001100110011001100110011","0001000000000000000000000000","0000001000010010000100100001","0000001110000011100000111000","0000011001000110010001100100","0000010001010100010101000101","0000001101010011010100110101","0000001001100010011000100110","0001000000000000000000000000","0000001001100010011000100110","0000011000010110000101100001","0000101000101010001010100010","0000011011100110111001101110","0000011000110110001101100011","0000011111000111110001111100","0000101110111011101110111011","0000111000111110001111100011","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111010101110101011101010","0000110101101101011011010110","0000110011001100110011001100","0000111010101110101011101010","0000100010011000100110001001","0000010100010101000101010001","0000111001001110010011100100","0000111110011111100111111001","0000111000101110001011100010","0000010100110101001101010011","0000010000110100001101000011","0000010100100101001001010010","0000010001010100010101000101","0000000001010000010100000101","0000100111001001110010011100","0000111001101110011011100110","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000110110111101101111011011","0000001101000011010000110100","0000000101010001010100010101","0000011000000110000001100000","0000100001101000011010000110","0000100001101000011010000110","0000100111101001111010011110","0000101011101010111010101110","0000100010101000101010001010","0000100100101001001010010010","0000001001000010010000100100","0000000111110001111100011111","0000101010101010101010101010","0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111011111110111111101","0000111100111111001111110011","0000111101011111010111110101","0000111111101111111011111110","0000111110101111101011111010","0000111101101111011011110110","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110011111100111111001","0000111101111111011111110111","0000111101011111010111110101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000110000111100001111000011","0000111000111110001111100011","0000100100011001000110010001","0000010111110101111101011111","0000101100011011000110110001","0000110001101100011011000110","0000011100110111001101110011","0000000110110001101100011011","0000000010000000100000001000","0000000101010001010100010101","0000010011000100110001001100","0000011110000111100001111000","0000100001011000010110000101","0000011100000111000001110000","0000010111010101110101011101","0000010010000100100001001000","0001000000000000000000000000","0000000000010000000100000001","0000000100110001001100010011","0000000100000001000000010000","0000011101000111010001110100","0000101001011010010110100101","0000101110101011101010111010","0000110010001100100011001000","0000111011111110111111101111","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000101101011011010110110101","0000100101001001010010010100","0000001111010011110100111101","0001000000000000000000000000","0000011010010110100101101001","0000001111000011110000111100","0000000011100000111000001110","0001000000000000000000000000","0000010111100101111001011110","0000110100111101001111010011","0000111010011110100111101001","0000111101001111010011110100","0000111100011111000111110001","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000100111111001111110011111","0000100000011000000110000001","0000011011000110110001101100","0000000101010001010100010101","0000001010010010100100101001","0000011101000111010001110100","0000000110100001101000011010","0000000110000001100000011000","0000001110110011101100111011","0000011101100111011001110110","0000011101010111010101110101","0000100111111001111110011111","0000101010101010101010101010","0000110110111101101111011011","0000111000101110001011100010","0000111010111110101111101011","0000111111111111111111111111","0000111111001111110011111100","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000100011111000111110001111","0000011000110110001101100011","0000101000111010001110100011","0000110101101101011011010110","0000101100111011001110110011","0000111110001111100011111000","0000111110001111100011111000","0000110111001101110011011100","0000111011001110110011101100","0000101100101011001010110010","0000110010101100101011001010","0000110101111101011111010111","0000110010001100100011001000","0000110101111101011111010111","0000111011101110111011101110","0000110110111101101111011011","0000101110011011100110111001","0000100110101001101010011010","0000011101000111010001110100","0000011101110111011101110111","0000100011111000111110001111","0000010000100100001001000010","0000000000100000001000000010","0000010110100101101001011010","0000010100000101000001010000","0000100011011000110110001101","0000111110111111101111111011","0000111010111110101111101011","0000111101111111011111110111","0000111111011111110111111101","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111001101110011011100110","0000101010111010101110101011","0000011110010111100101111001","0000100011111000111110001111","0000011101010111010101110101","0001000000000000000000000000","0000001011000010110000101100","0000010011010100110101001101","0000011001110110011101100111","0000011100010111000101110001","0000100001011000010110000101","0000011110000111100001111000","0000100010111000101110001011","0000100101001001010010010100","0000011101000111010001110100","0000010111100101111001011110","0000000011100000111000001110","0000010100010101000101010001","0000011001000110010001100100","0000100000111000001110000011","0000011100000111000001110000","0000100100101001001010010010","0000101000001010000010100000","0000100101011001010110010101","0000101100111011001110110011","0000100101101001011010010110","0000110100101101001011010010","0000110011011100110111001101","0000010111110101111101011111","0000010001110100011101000111","0000100101111001011110010111","0000111011001110110011101100","0000111110111111101111111011","0000111111111111111111111111","0000100000001000000010000000","0000001011110010111100101111","0000010001110100011101000111","0000011110000111100001111000","0001000000000000000000000000","0000011110000111100001111000","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101011111010111110101","0000111111111111111111111111","0000111011011110110111101101","0000100100101001001010010010","0000000011010000110100001101","0000000110010001100100011001","0000011011000110110001101100","0000100011001000110010001100","0000101111101011111010111110","0000111100011111000111110001","0000111101111111011111110111","0000110111111101111111011111","0000011001010110010101100101","0000001010110010101100101011","0000010100100101001001010010","0000100101001001010010010100","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111011001110110011101100","0000111101001111010011110100","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111001111110011111100111","0000110111001101110011011100","0000110010101100101011001010","0000011111000111110001111100","0000100011001000110010001100","0000100110111001101110011011","0000011101000111010001110100","0000000100010001000100010001","0000000101100001011000010110","0000100101101001011010010110","0000100110111001101110011011","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111001111110011111100111","0000111111111111111111111111","0000111000111110001111100011","0000100101011001010110010101","0000010000100100001001000010","0000010011000100110001001100","0000010010100100101001001010","0000011001010110010101100101","0000101011011010110110101101","0000111010011110100111101001","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000100110101001101010011010","0000010100100101001001010010","0000001001000010010000100100","0000000010110000101100001011","0000011000000110000001100000","0000010111100101111001011110","0000010011010100110101001101","0000000000100000001000000010","0000010101000101010001010100","0000100100111001001110010011","0000110110101101101011011010","0000111100101111001011110010","0000111100011111000111110001","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000100101111001011110010111","0000011100010111000101110001","0000011010000110100001101000","0000000110000001100000011000","0000001001100010011000100110","0000001011110010111100101111","0000011100100111001001110010","0000011111000111110001111100","0000010100100101001001010010","0000010000110100001101000011","0000011111110111111101111111","0000110010001100100011001000","0000111001001110010011100100","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000110110111101101111011011","0000100110101001101010011010","0000101111011011110110111101","0000110100011101000111010001","0000111010101110101011101010","0000111110011111100111111001","0000111110111111101111111011","0000111101001111010011110100","0000111010111110101111101011","0000111111111111111111111111","0000111111001111110011111100","0000110101001101010011010100","0000110110111101101111011011","0000110011111100111111001111","0000101100011011000110110001","0000100000001000000010000000","0000011001100110011001100110","0000011101010111010101110101","0000011110000111100001111000","0000101001101010011010100110","0000100111011001110110011101","0000001011000010110000101100","0000010010100100101001001010","0000011011110110111101101111","0000001100010011000100110001","0000110011001100110011001100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100001111000011110000","0000111011111110111111101111","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111011111110111111101111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100011101000111010001","0000100001111000011110000111","0000100101101001011010010110","0000101100111011001110110011","0000100010001000100010001000","0000001001110010011100100111","0000011001110110011101100111","0000001100110011001100110011","0000001011000010110000101100","0000001100010011000100110001","0000001100100011001000110010","0000100100011001000110010001","0000110011001100110011001100","0000110001011100010111000101","0000111011001110110011101100","0000111011001110110011101100","0000110110011101100111011001","0000011111000111110001111100","0000000011110000111100001111","0000000100110001001100010011","0000011011010110110101101101","0000011101000111010001110100","0000011111100111111001111110","0000100111011001110110011101","0000100001101000011010000110","0000101110111011101110111011","0000101101111011011110110111","0000100001001000010010000100","0001000000000000000000000000","0000100001001000010010000100","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000101010111010101110101011","0000100000001000000010000000","0000010110100101101001011010","0000010101110101011101010111","0000000110110001101100011011","0000010100000101000001010000","0000111101101111011011110110","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111111011111110111111101","0000111001011110010111100101","0000001110010011100100111001","0000000110000001100000011000","0000001000000010000000100000","0000011111010111110101111101","0000101000111010001110100011","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000101001011010010110100101","0000001001000010010000100100","0000001100010011000100110001","0000011110000111100001111000","0000110111101101111011011110","0000111011011110110111101101","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111101011111010111110101","0000111111001111110011111100","0000111110101111101011111010","0000111101001111010011110100","0000111100101111001011110010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111101101111011011110110","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111000001110000011100000","0000010111010101110101011101","0000100101001001010010010100","0000100111011001110110011101","0000100010111000101110001011","0000001011100010111000101110","0000011000110110001101100011","0000011010110110101101101011","0000110000001100000011000000","0000101111101011111010111110","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000110011101100111011001110","0000100000001000000010000000","0000011111010111110101111101","0000011100110111001101110011","0000011111000111110001111100","0000100101011001010110010101","0000101001111010011110100111","0000110010111100101111001011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111001101110011011100110","0000010110110101101101011011","0000000111110001111100011111","0000000100110001001100010011","0000001110110011101100111011","0000010011110100111101001111","0000010010010100100101001001","0000011101000111010001110100","0000010100010101000101010001","0000000100010001000100010001","0000100111011001110110011101","0000110010101100101011001010","0000111000101110001011100010","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111100111111001111110011","0000100011011000110110001101","0000101110011011100110111001","0000000100100001001000010010","0000000011110000111100001111","0000000101010001010100010101","0000010011010100110101001101","0000011000010110000101100001","0000100000101000001010000010","0000011000110110001101100011","0000101110001011100010111000","0000110011001100110011001100","0000110101001101010011010100","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111011111110111111101111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000110111101101111011011110","0000111000001110000011100000","0000110110001101100011011000","0000111111111111111111111111","0000111010011110100111101001","0000111001101110011011100110","0000111001111110011111100111","0000111101111111011111110111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000110011101100111011001110","0000100101001001010010010100","0000100000101000001010000010","0000100110101001101010011010","0000110010111100101111001011","0000110110011101100111011001","0000100101001001010010010100","0000010011100100111001001110","0000000011000000110000001100","0000011110110111101101111011","0000101010111010101110101011","0000010000110100001101000011","0000110010001100100011001000","0000111000001110000011100000","0000111010101110101011101010","0000111101011111010111110101","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111111101111111011111110","0000111111011111110111111101","0000111110011111100111111001","0000111101001111010011110100","0000110111001101110011011100","0000100110011001100110011001","0000010100010101000101010001","0000100101101001011010010110","0000111110101111101011111010","0000000111000001110000011100","0000011010100110101001101010","0000001111100011111000111110","0000011001100110011001100110","0000011000000110000001100000","0000011001100110011001100110","0000100010001000100010001000","0000011110100111101001111010","0000101011101010111010101110","0000111110001111100011111000","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000100001011000010110000101","0000000001000000010000000100","0000001100010011000100110001","0000010111110101111101011111","0000010100100101001001010010","0000100010001000100010001000","0000100100111001001110010011","0000100010011000100110001001","0000000010100000101000001010","0000100101001001010010010100","0000111111001111110011111100","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000101111101011111010111110","0000011011010110110101101101","0000001000010010000100100001","0000010001100100011001000110","0000011110010111100101111001","0001000000000000000000000000","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101111111011111110111","0000111111111111111111111111","0000110000011100000111000001","0000001011110010111100101111","0001000000000000000000000000","0000010111110101111101011111","0000011010110110101101101011","0000110011111100111111001111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000110011101100111011001110","0000001110010011100100111001","0000100010101000101010001010","0000001111010011110100111101","0000110001011100010111000101","0000111100111111001111110011","0000111111011111110111111101","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000110100001101000011010000","0000101110111011101110111011","0000101110001011100010111000","0000101111011011110110111101","0000111101111111011111110111","0000111110001111100011111000","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111111111111111111111111","0000111101001111010011110100","0000100010111000101110001011","0000100010011000100110001001","0000100001001000010010000100","0000110001001100010011000100","0000001010000010100000101000","0000100110001001100010011000","0000011101100111011001110110","0000101010111010101110101011","0000111010111110101111101011","0000111010111110101111101011","0000111110011111100111111001","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000101101011011010110110101","0000100011001000110010001100","0000101101011011010110110101","0000111011111110111111101111","0000111111011111110111111101","0000111000101110001011100010","0000110001011100010111000101","0000111000011110000111100001","0000111011101110111011101110","0000110100001101000011010000","0000010111010101110101011101","0000010000010100000101000001","0000000001110000011100000111","0000010100100101001001010010","0000011010000110100001101000","0000100100011001000110010001","0000011101100111011001110110","0000011011000110110001101100","0001000000000000000000000000","0000010001000100010001000100","0000110010011100100111001001","0000111010011110100111101001","0000111100001111000011110000","0000111110111111101111111011","0000111101001111010011110100","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110111111101111111011","0000111011101110111011101110","0000100001101000011010000110","0000010000010100000101000001","0000000001010000010100000101","0000001100000011000000110000","0000000111110001111100011111","0000010100100101001001010010","0000100000011000000110000001","0000100011001000110010001100","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111100111111001111110011","0000111111001111110011111100","0000111101001111010011110100","0000111111011111110111111101","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111011011110110111101101","0000111111011111110111111101","0000111111111111111111111111","0000110110101101101011011010","0000111010001110100011101000","0000111110011111100111111001","0000110100001101000011010000","0000111111111111111111111111","0000111100111111001111110011","0000111110001111100011111000","0000110010011100100111001001","0000110111011101110111011101","0000101010111010101110101011","0000101011001010110010101100","0000101101001011010010110100","0000101000001010000010100000","0000011010010110100101101001","0000011110100111101001111010","0000101011101010111010101110","0000101010111010101110101011","0000100001011000010110000101","0000010101110101011101010111","0000000001110000011100000111","0000000011010000110100001101","0000011100000111000001110000","0000011110100111101001111010","0000101011011010110110101101","0000001110000011100000111000","0000001101000011010000110100","0000110111101101111011011110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111011011110110111101101","0000101101001011010010110100","0000011111100111111001111110","0000101110011011100110111001","0000010111110101111101011111","0000000011100000111000001110","0001000000000000000000000000","0000100100011001000110010001","0000101010011010100110101001","0000110011101100111011001110","0000110100111101001111010011","0000101001011010010110100101","0000100100011001000110010001","0000100000011000000110000001","0000110011001100110011001100","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000100000111000001110000011","0000001001010010010100100101","0000000010100000101000001010","0001000000000000000000000000","0001000000000000000000000000","0000000010110000101100001011","0000101011101010111010101110","0000111101001111010011110100","0000111110001111100011111000","0000111111011111110111111101","0000111100101111001011110010","0000111110101111101011111010","0000111111111111111111111111","0000110010001100100011001000","0000100101011001010110010101","0000010011000100110001001100","0000010111100101111001011110","0000011101000111010001110100","0000000010110000101100001011","0000101010111010101110101011","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110101111101011111010","0000111101111111011111110111","0000110111011101110111011101","0001000000000000000000000000","0000000101110001011100010111","0000011110010111100101111001","0000011110110111101101111011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111100011111000111110001","0000101100001011000010110000","0000100010101000101010001010","0000011011100110111001101110","0000001111110011111100111111","0000101000101010001010100010","0000111010011110100111101001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000110011011100110111001101","0000101010111010101110101011","0000100100101001001010010010","0000110010001100100011001000","0000110010101100101011001010","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111101111111011111110","0000111000111110001111100011","0000100101111001011110010111","0000110101101101011011010110","0000111111111111111111111111","0000111001111110011111100111","0000111111111111111111111111","0000111111001111110011111100","0000111010101110101011101010","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000110101111101011111010111","0000011111010111110101111101","0000100000111000001110000011","0000101110011011100110111001","0000010010100100101001001010","0000101011011010110110101101","0000101000111010001110100011","0000101100111011001110110011","0000110111111101111111011111","0000111100101111001011110010","0000111110001111100011111000","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111000011110000111100001","0000100010111000101110001011","0000110101101101011011010110","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111011011110110111101101","0000111111001111110011111100","0000100001101000011010000110","0000010000110100001101000011","0000001010010010100100101001","0001000000000000000000000000","0000011011100110111001101110","0000010111010101110101011101","0000010111100101111001011110","0000010110010101100101011001","0000010100000101000001010000","0000001100100011001000110010","0001000000000000000000000000","0000100010011000100110001001","0000100111001001110010011100","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000101010111010101110101011","0000011001100110011001100110","0000010001010100010101000101","0000001101110011011100110111","0000000110110001101100011011","0000001100100011001000110010","0000011011110110111101101111","0000101111001011110010111100","0000111100111111001111110011","0000111010101110101011101010","0000111100001111000011110000","0000111110101111101011111010","0000111111001111110011111100","0000111110011111100111111001","0000111111001111110011111100","0000111111011111110111111101","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000110110111101101111011011","0000111101001111010011110100","0000110011101100111011001110","0000110101101101011011010110","0000111011011110110111101101","0000111011111110111111101111","0000101111001011110010111100","0000011111100111111001111110","0000100111011001110110011101","0000011011000110110001101100","0000011000100110001001100010","0000010000110100001101000011","0000010100000101000001010000","0000011001000110010001100100","0000010011000100110001001100","0000010110100101101001011010","0000000100010001000100010001","0000001000100010001000100010","0000001110110011101100111011","0000010101000101010001010100","0000010010010100100101001001","0000010110100101101001011010","0000010011000100110001001100","0000100010111000101110001011","0000101001011010010110100101","0000110001111100011111000111","0000111011001110110011101100","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111011011110110111101101","0000111110101111101011111010","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000110111101101111011011110","0000110000101100001011000010","0000101011111010111110101111","0000110000101100001011000010","0000100001001000010010000100","0001000000000000000000000000","0000011111110111111101111111","0000110110101101101011011010","0000101111101011111010111110","0000101101111011011110110111","0000110110101101101011011010","0000110101011101010111010101","0000111110101111101011111010","0000110111101101111011011110","0000101010101010101010101010","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111011011110110111101101","0000110100011101000111010001","0000111100011111000111110001","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111110101111101011111010","0000111101001111010011110100","0000111100111111001111110011","0000111011111110111111101111","0000110000111100001111000011","0000100011111000111110001111","0000011001100110011001100110","0000100111101001111010011110","0000010110000101100001011000","0000000100000001000000010000","0000101111011011110110111101","0000111001001110010011100100","0000111111101111111011111110","0000111111101111111011111110",
		"0000111011011110110111101101","0000111111111111111111111111","0000110001001100010011000100","0001000000000000000000000000","0000001011100010111000101110","0000011000010110000101100001","0000101110001011100010111000","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111000101110001011100010","0000111010011110100111101001","0000111111111111111111111111","0000101001111010011110100111","0000001010100010101000101010","0000000110000001100000011000","0000010110000101100001011000","0000110110111101101111011011","0000111111111111111111111111","0000111011011110110111101101","0000111010011110100111101001","0000111111111111111111111111","0000111101101111011011110110","0000110000011100000111000001","0000101101011011010110110101","0000010110010101100101011001","0000100010011000100110001001","0000100010101000101010001010","0000111001111110011111100111","0000111111111111111111111111","0000111001001110010011100100","0000110101111101011111010111","0000110111111101111111011111","0000101001001010010010100100","0000111000011110000111100001","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111111111111111111111111","0000111001011110010111100101","0000111100001111000011110000","0000111111111111111111111111","0000111111011111110111111101","0000101011111010111110101111","0000100111111001111110011111","0000100000101000001010000010","0000101011101010111010101110","0000001110010011100100111001","0000101000111010001110100011","0000110010111100101111001011","0000111011011110110111101101","0000110111101101111011011110","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000110001001100010011000100","0000110100001101000011010000","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000110111001101110011011100","0000100000001000000010000000","0000011001000110010001100100","0000001011010010110100101101","0000000000110000001100000011","0000010110000101100001011000","0000100011101000111010001110","0000101000111010001110100011","0000100001101000011010000110","0000011100100111001001110010","0000010010000100100001001000","0000000000010000000100000001","0000011011110110111101101111","0000100000111000001110000011","0000110011001100110011001100","0000111111011111110111111101","0000111100001111000011110000","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000011110110111101101111011","0000010101000101010001010100","0000010010000100100001001000","0000001110010011100100111001","0001000000000000000000000000","0000011010010110100101101001","0000100011001000110010001100","0000111000101110001011100010","0000101101111011011110110111","0000111011001110110011101100","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111000111110001111100011","0000110001101100011011000110","0000101100011011000110110001","0000100000111000001110000011","0000011110100111101001111010","0000011110000111100001111000","0000011110010111100101111001","0000011001010110010101100101","0000100100011001000110010001","0000100000001000000010000000","0000011110000111100001111000","0000011010100110101001101010","0000010011000100110001001100","0000001101110011011100110111","0000001010000010100000101000","0000010100010101000101010001","0000001110110011101100111011","0000001001010010010100100101","0000010000100100001001000010","0000100000001000000010000000","0000011100010111000101110001","0000011010100110101001101010","0000011010000110100001101000","0000011110100111101001111010","0000011101000111010001110100","0000011110000111100001111000","0000100101011001010110010101","0000101001011010010110100101","0000110001101100011011000110","0000110110111101101111011011","0000110000011100000111000001","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000110111001101110011011100","0000110000111100001111000011","0000101110111011101110111011","0000101011001010110010101100","0000100001001000010010000100","0000000010010000100100001001","0000100011101000111010001110","0000101110011011100110111001","0000100011101000111010001110","0000101100101011001010110010","0000101011101010111010101110","0000111101011111010111110101","0000111101011111010111110101","0000111010011110100111101001","0000111011001110110011101100","0000110010011100100111001001","0000111110011111100111111001","0000111111111111111111111111","0000111011111110111111101111","0000111101111111011111110111","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000111100111111001111110011","0000111111101111111011111110","0000111110001111100011111000","0000111100001111000011110000","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000110000101100001011000010","0000011110110111101101111011","0000011000110110001101100011","0000101100111011001110110011","0001000000000000000000000000","0000010100000101000001010000","0000110101001101010011010100","0000111011001110110011101100","0000111111101111111011111110","0000111111101111111011111110",
		"0000111011101110111011101110","0000111111111111111111111111","0000101010101010101010101010","0000000010100000101000001010","0000001110110011101100111011","0000010111100101111001011110","0000111001001110010011100100","0000111101111111011111110111","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111001111110011111100111","0000101111001011110010111100","0000101100111011001110110011","0000100001011000010110000101","0000001001000010010000100100","0000000000010000000100000001","0000010101010101010101010101","0000101011001010110010101100","0000110000111100001111000011","0000101100011011000110110001","0000100001011000010110000101","0000010100100101001001010010","0000010000110100001101000011","0000001011010010110100101101","0000010011010100110101001101","0000000111010001110100011101","0001000000000000000000000000","0000000100110001001100010011","0000010100110101001101010011","0000110010011100100111001001","0000110111011101110111011101","0000101100001011000010110000","0000110000001100000011000000","0000101001111010011110100111","0000110010001100100011001000","0000111110011111100111111001","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000101101101011011010110110","0000100111001001110010011100","0000101111101011111010111110","0000010101000101010001010100","0000010111100101111001011110","0000101010011010100110101001","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111110101111101011111010","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000110011001100110011001100","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000110100001101000011010000","0000100011001000110010001100","0000011110010111100101111001","0000001101010011010100110101","0000001000110010001100100011","0000010110110101101101011011","0000100000101000001010000010","0000100111111001111110011111","0000100010011000100110001001","0000100011111000111110001111","0000011111100111111001111110","0000001110010011100100111001","0001000000000000000000000000","0000011001010110010101100101","0000100110111001101110011011","0000101110101011101010111010","0000111110001111100011111000","0000111111111111111111111111","0000111010101110101011101010","0000110011011100110111001101","0000100011011000110110001101","0000010000100100001001000010","0000001111000011110000111100","0000010011100100111001001110","0000010110000101100001011000","0001000000000000000000000000","0000011000000110000001100000","0000101000101010001010100010","0000110100101101001011010010","0000110000101100001011000010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111001001110010011100100","0000111100011111000111110001","0000111001101110011011100110","0000110101001101010011010100","0000110011111100111111001111","0000110001101100011011000110","0000100111011001110110011101","0000011010010110100101101001","0000010110000101100001011000","0000011010100110101001101010","0000100101011001010110010101","0000101011011010110110101101","0000011111110111111101111111","0000011101010111010101110101","0000001110110011101100111011","0000001111000011110000111100","0000001011010010110100101101","0000010000110100001101000011","0000011000100110001001100010","0000010110010101100101011001","0000100100001001000010010000","0000011100000111000001110000","0000100001111000011110000111","0000011111110111111101111111","0000011101110111011101110111","0000011010110110101101101011","0000010001100100011001000110","0000010011000100110001001100","0000011101110111011101110111","0000011110100111101001111010","0000100100001001000010010000","0000101011101010111010101110","0000101001011010010110100101","0000101011111010111110101111","0000100101101001011010010110","0000101010101010101010101010","0000100110101001101010011010","0000111000101110001011100010","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000110111001101110011011100","0000110001011100010111000101","0000110011101100111011001110","0000110001111100011111000111","0000100010111000101110001011","0000000101000001010000010100","0000011111010111110101111101","0000011010110110101101101011","0000100011111000111110001111","0000100101111001011110010111","0000110100011101000111010001","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000110111111101111111011111","0000110111111101111111011111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111110111111101111111011","0000111011101110111011101110","0000111010111110101111101011","0000111111111111111111111111","0000110110001101100011011000","0000010111110101111101011111","0000011110000111100001111000","0000101100111011001110110011","0000000011010000110100001101","0000011010010110100101101001","0000110010111100101111001011","0000111010101110101011101010","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111111111111111111111","0000111101111111011111110111","0000101001001010010010100100","0000000110110001101100011011","0000001011100010111000101110","0000011110000111100001111000","0000111001001110010011100100","0000111110011111100111111001","0000111110001111100011111000","0000111101001111010011110100","0000111110001111100011111000","0000111010001110100011101000","0000101110111011101110111011","0000100111001001110010011100","0000100101101001011010010110","0000100100101001001010010010","0000010101100101011001010110","0000011100100111001001110010","0000011001010110010101100101","0000000100110001001100010011","0000000011010000110100001101","0000010101110101011101010111","0000011011110110111101101111","0000011010010110100101101001","0000011011110110111101101111","0000100010011000100110001001","0000100111011001110110011101","0000100111101001111010011110","0000100000011000000110000001","0000010111100101111001011110","0000000000100000001000000010","0000011111110111111101111111","0000100111101001111010011110","0000101011101010111010101110","0000110000111100001111000011","0000100100001001000010010000","0000111000001110000011100000","0000111111111111111111111111","0000111101011111010111110101","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111101011111010111110101","0000110100111101001111010011","0000100100001001000010010000","0000110010011100100111001001","0001000000000000000000000000","0000100001101000011010000110","0000110011001100110011001100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000110101101101011011010110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000110110001101100011011000","0000111101001111010011110100","0000111110101111101011111010","0000111111001111110011111100","0000111111101111111011111110","0000110011001100110011001100","0000011101000111010001110100","0000011000110110001101100011","0000000101000001010000010100","0000001011110010111100101111","0000010111110101111101011111","0000011011110110111101101111","0000100010101000101010001010","0000110010011100100111001001","0000111010001110100011101000","0000101000011010000110100001","0000010001110100011101000111","0000010111000101110001011100","0000010100010101000101010001","0000001111110011111100111111","0000011110100111101001111010","0000101000101010001010100010","0000101111101011111010111110","0000110011111100111111001111","0000101011111010111110101111","0000010011000100110001001100","0000001010000010100000101000","0000011000000110000001100000","0000010001000100010001000100","0000011101010111010101110101","0000000000110000001100000011","0000010110100101101001011010","0000101001111010011110100111","0000101001011010010110100101","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111010101110101011101010","0000111111111111111111111111","0000111100001111000011110000","0000101011001010110010101100","0000101110011011100110111001","0000110101001101010011010100","0000110011111100111111001111","0000110001001100010011000100","0000101101101011011010110110","0000101000101010001010100010","0000100010011000100110001001","0000010110110101101101011011","0000011110000111100001111000","0000100001011000010110000101","0000011010100110101001101010","0000011000000110000001100000","0000010111010101110101011101","0000100001101000011010000110","0000100001001000010010000100","0000100010111000101110001011","0000100111101001111010011110","0000011111010111110101111101","0000001000110010001100100011","0000001111010011110100111101","0000010100000101000001010000","0000001001000010010000100100","0000001100100011001000110010","0000001110110011101100111011","0000001110100011101000111010","0000000110100001101000011010","0001000000000000000000000000","0000000100100001001000010010","0000001001110010011100100111","0000010101100101011001010110","0000011001000110010001100100","0000011111010111110101111101","0000100001111000011110000111","0000100010011000100110001001","0000100000111000001110000011","0000100001011000010110000101","0000111000001110000011100000","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000110111111101111111011111","0000110001111100011111000111","0000111000111110001111100011","0000110100111101001111010011","0000100010001000100010001000","0001000000000000000000000000","0000010101100101011001010110","0000001110000011100000111000","0000011100000111000001110000","0000100011001000110010001100","0000111110111111101111111011","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111001011110010111100101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111011111110111111101","0000111010001110100011101000","0000111111001111110011111100","0000111010001110100011101000","0000111111101111111011111110","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110100001101000011010000","0000111000101110001011100010","0000101101001011010010110100","0000100100011001000110010001","0000110100111101001111010011","0000101101011011010110110101","0000010110000101100001011000","0000001001100010011000100110","0000100110101001101010011010","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111111111111111111111","0000111110001111100011111000","0000101101001011010010110100","0000000100110001001100010011","0000000111100001111000011110","0000100010001000100010001000","0000111010011110100111101001","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111001111110011111100","0000101100101011001010110010","0000011110100111101001111010","0000100100101001001010010010","0000011000000110000001100000","0000010010110100101101001011","0000011000100110001001100010","0000011110100111101001111010","0000100101111001011110010111","0000101110001011100010111000","0000110001101100011011000110","0000111000111110001111100011","0000111011001110110011101100","0000111001101110011011100110","0000111110101111101011111010","0000111111111111111111111111","0000110001111100011111000111","0000101000101010001010100010","0000100010011000100110001001","0001000000000000000000000000","0000100011001000110010001100","0000100000101000001010000010","0000101010101010101010101010","0000110011001100110011001100","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111000111110001111100011","0000110010101100101011001010","0000101000101010001010100010","0000011111110111111101111111","0000000010010000100100001001","0000011110100111101001111010","0000111000111110001111100011","0000111111111111111111111111","0000110110011101100111011001","0000111110111111101111111011","0000101110101011101010111010","0000111101011111010111110101","0000111100001111000011110000","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000111100111111001111110011","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000110110101101101011011010","0000101000111010001110100011","0000010101010101010101010101","0000100001101000011010000110","0000000010010000100100001001","0000010100010101000101010001","0000001110100011101000111010","0000011111110111111101111111","0000110000011100000111000001","0000110111001101110011011100","0000111010111110101111101011","0000111010001110100011101000","0000110110111101101111011011","0000011101100111011001110110","0000011001010110010101100101","0000010110100101101001011010","0000000101100001011000010110","0000010000110100001101000011","0000010101110101011101010111","0000010011100100111001001110","0000010000010100000101000001","0000001111100011111000111110","0000011000110110001101100011","0000100110101001101010011010","0000001011010010110100101101","0000011001110110011101100111","0000000000110000001100000011","0000100010111000101110001011","0000101000001010000010100000","0000101011101010111010101110","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000110011001100110011001100","0000101110101011101010111010","0000111010011110100111101001","0000110110111101101111011011","0000101111111011111110111111","0000101000111010001110100011","0000110100001101000011010000","0000111100111111001111110011","0000111001111110011111100111","0000111000111110001111100011","0000110011111100111111001111","0000101101001011010010110100","0000100010101000101010001010","0000011000110110001101100011","0000011111110111111101111111","0000100100101001001010010010","0000101011011010110110101101","0000011110110111101101111011","0000010010010100100101001001","0000010111010101110101011101","0000001100010011000100110001","0000001111000011110000111100","0000100100101001001010010010","0000101011111010111110101111","0000110110111101101111011011","0000110101111101011111010111","0000111000101110001011100010","0000111011111110111111101111","0000101110011011100110111001","0000011001110110011101100111","0000100001001000010010000100","0000011101110111011101110111","0000001110110011101100111011","0000000111100001111000011110","0001000000000000000000000000","0000010010010100100101001001","0000011101110111011101110111","0000100011111000111110001111","0000100110101001101010011010","0000100001011000010110000101","0000110100101101001011010010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111001111110011111100111","0000110010001100100011001000","0000111101001111010011110100","0000110110101101101011011010","0000100110111001101110011011","0000000001010000010100000101","0000100011001000110010001100","0000010011110100111101001111","0000010000010100000101000001","0000110000001100000011000000","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111100011111000111110001","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111011111110111111101111","0000110100111101001111010011","0000111111111111111111111111","0000110001111100011111000111","0000111111111111111111111111","0000111010101110101011101010","0000111011001110110011101100","0000111111111111111111111111","0000111100111111001111110011","0000111101001111010011110100","0000111111111111111111111111","0000101101101011011010110110","0000110111101101111011011110","0000100110011001100110011001","0000111011011110110111101101","0000111111001111110011111100","0000100110011001100110011001","0000011011010110110101101101","0000000000100000001000000010","0000100010011000100110001001","0000111110101111101011111010","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111001111110011111100","0000111111111111111111111111","0000110000111100001111000011","0001000000000000000000000000","0000000110010001100100011001","0000011111100111111001111110","0000111110111111101111111011","0000110001101100011011000110","0000111011001110110011101100","0000111011011110110111101101","0000111111101111111011111110","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000101111011011110110111101","0000101011001010110010101100","0000100101001001010010010100","0000101000001010000010100000","0000101100011011000110110001","0000101100111011001110110011","0000101110011011100110111001","0000110000111100001111000011","0000110100111101001111010011","0000111010101110101011101010","0000111101111111011111110111","0000111101011111010111110101","0000111110011111100111111001","0000111111111111111111111111","0000110101011101010111010101","0000111000001110000011100000","0000101101101011011010110110","0000000000010000000100000001","0000100010011000100110001001","0000100010101000101010001010","0000101101001011010010110100","0000101100111011001110110011","0000111111001111110011111100","0000111110001111100011111000","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111100001111000011110000","0000110001101100011011000110","0000101001001010010010100100","0000010111010101110101011101","0000010000100100001001000010","0000011101010111010101110101","0000111001101110011011100110","0000110110111101101111011011","0000111111111111111111111111","0000100111111001111110011111","0000111100001111000011110000","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000100011001000110010001100","0000011110110111101101111011","0000001011000010110000101100","0000000111000001110000011100","0000010010100100101001001010","0000100001111000011110000111","0000111100001111000011110000","0000111100001111000011110000","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000100011101000111010001110","0000101111011011110110111101","0000101000001010000010100000","0000011100100111001001110010","0000010100100101001001010010","0000010011110100111101001111","0000010100010101000101010001","0000001111110011111100111111","0000010010000100100001001000","0000100001001000010010000100","0000001000110010001100100011","0000010010010100100101001001","0000001001110010011100100111","0000100001011000010110000101","0000100011011000110110001101","0000110010111100101111001011","0000111111101111111011111110","0000111110001111100011111000","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000110101111101011111010111","0000111010001110100011101000","0000111111101111111011111110","0000111011111110111111101111","0000111001001110010011100100","0000111111011111110111111101","0000111101001111010011110100","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000110010011100100111001001","0000100110111001101110011011","0000010111000101110001011100","0000000111110001111100011111","0000011001000110010001100100","0000011100110111001101110011","0000100010111000101110001011","0000010110010101100101011001","0000001110010011100100111001","0000000110000001100000011000","0000011111100111111001111110","0000100111111001111110011111","0000110000101100001011000010","0000101110101011101010111010","0000101110011011100110111001","0000111100101111001011110010","0000111101011111010111110101","0000111111111111111111111111","0000111010001110100011101000","0000100111101001111010011110","0000101000001010000010100000","0000110010001100100011001000","0000101001001010010010100100","0000110000001100000011000000","0000011111010111110101111101","0000001101100011011000110110","0000010011000100110001001100","0000001010100010101000101010","0000001001010010010100100101","0000101101011011010110110101","0000011111110111111101111111","0000110000011100000111000001","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111111001111110011111100","0000111100101111001011110010","0000110010011100100111001001","0000111111101111111011111110","0000110111101101111011011110","0000100100001001000010010000","0000000001010000010100000101","0000110001001100010011000100","0000000111010001110100011101","0000001111000011110000111100","0000101010101010101010101010","0000111101101111011011110110","0000111101111111011111110111","0000111111101111111011111110","0000111110101111101011111010","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111011001110110011101100","0000111110001111100011111000","0000111111111111111111111111","0000111011011110110111101101","0000111000011110000111100001","0000110001111100011111000111","0000111111111111111111111111","0000101111011011110110111101","0000111111011111110111111101","0000110101101101011011010110","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111100101111001011110010","0000110101111101011111010111","0000100110101001101010011010","0000101101101011011010110110","0000110001001100010011000100","0000111111111111111111111111","0000111001101110011011100110","0000011101110111011101110111","0000011111110111111101111111","0001000000000000000000000000","0000100111001001110010011100","0000111100111111001111110011","0000111111101111111011111110","0000111111101111111011111110",
		"0000111110111111101111111011","0000111111111111111111111111","0000110000011100000111000001","0001000000000000000000000000","0000000101010001010100010101","0000011101100111011001110110","0000111011001110110011101100","0000110001001100010011000100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111100111111001111110011","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111100011111000111110001","0000111010101110101011101010","0000111111111111111111111111","0000011111110111111101111111","0000001111110011111100111111","0000100110011001100110011001","0000110100001101000011010000","0000110101001101010011010100","0000110000001100000011000000","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111001001110010011100100","0000100110111001101110011011","0000010000010100000101000001","0000100001001000010010000100","0000100011111000111110001111","0000110000011100000111000001","0000110001011100010111000101","0000111000011110000111100001","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111011101110111011101110","0000111101111111011111110111","0000111101111111011111110111","0000111110011111100111111001","0000101011001010110010101100","0000011011010110110101101101","0000001110100011101000111010","0000001111000011110000111100","0000100001111000011110000111","0000101111111011111110111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000110110011101100111011001","0000100101101001011010010110","0000101010111010101110101011","0000101010101010101010101010","0000100000101000001010000010","0000100000001000000010000000","0000011011110110111101101111","0000010010100100101001001010","0000011100010111000101110001","0000001000000010000000100000","0000010000000100000001000000","0000010011100100111001001110","0000011000110110001101100011","0000100000101000001010000010","0000101110001011100010111000","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111010011110100111101001","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000110101111101011111010111","0000100110111001101110011011","0000001011110010111100101111","0000010000100100001001000010","0000010111010101110101011101","0000011001010110010101100101","0000010001100100011001000110","0000001010010010100100101001","0000001010010010100100101001","0000011111100111111001111110","0000101010111010101110101011","0000101010001010100010101000","0000111011001110110011101100","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111101101111011011110110","0000111100111111001111110011","0000101100101011001010110010","0000100100011001000110010001","0000101111101011111010111110","0000110000011100000111000001","0000111110111111101111111011","0000101111011011110110111101","0000100111011001110110011101","0000010000000100000001000000","0000010111010101110101011101","0000010001100100011001000110","0000010001100100011001000110","0000010001100100011001000110","0000100100001001000010010000","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000110010011100100111001001","0000111111111111111111111111","0000111101011111010111110101","0000100111101001111010011110","0000000010100000101000001010","0000110000101100001011000010","0000000100100001001000010010","0000011100100111001001110010","0000100001101000011010000110","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111010011110100111101001","0000111110011111100111111001","0000111111111111111111111111","0000111001011110010111100101","0000110100101101001011010010","0000101111001011110010111100","0000110101101101011011010110","0000110000011100000111000001","0000110111001101110011011100","0000101111001011110010111100","0000111010111110101111101011","0000111101011111010111110101","0000111111111111111111111111","0000110111101101111011011110","0000100101111001011110010111","0000010100010101000101010001","0000100100011001000110010001","0000111001111110011111100111","0000111001011110010111100101","0000111011001110110011101100","0000100101101001011010010110","0000101011001010110010101100","0001000000000000000000000000","0000100100011001000110010001","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111111111111111111111","0000111011011110110111101101","0000101101101011011010110110","0000000001000000010000000100","0000000011100000111000001110","0000011111000111110001111100","0000110001101100011011000110","0000110101111101011111010111","0000110101011101010111010101","0000110111111101111111011111","0000111011111110111111101111","0000111111101111111011111110","0000111111101111111011111110","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111011001110110011101100","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111100001111000011110000","0000000011000000110000001100","0000100001011000010110000101","0000101010011010100110101001","0000110001111100011111000111","0000111000101110001011100010","0000111110001111100011111000","0000111110101111101011111010","0000111110011111100111111001","0000111110011111100111111001","0000111011101110111011101110","0000111111011111110111111101","0000101001101010011010100110","0001000000000000000000000000","0000110010001100100011001000","0000100111001001110010011100","0000100111001001110010011100","0000101110101011101010111010","0000100111011001110110011101","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111011111110111111101","0000111100111111001111110011","0000111000101110001011100010","0000111000101110001011100010","0000111000101110001011100010","0000111000101110001011100010","0000111000101110001011100010","0000111000101110001011100010","0000111000101110001011100010","0000111000101110001011100010","0000111011011110110111101101","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111000101110001011100010","0000111011001110110011101100","0000111000101110001011100010","0000110111011101110111011101","0000100111001001110010011100","0000011001010110010101100101","0000001000100010001000100010","0000101000011010000110100001","0000011011010110110101101101","0000111011001110110011101100","0000101111111011111110111111","0000101011101010111010101110","0000101101011011010110110101","0000110001001100010011000100","0000110011011100110111001101","0000110000101100001011000010","0000110000101100001011000010","0000110101111101011111010111","0000111111001111110011111100","0000111111101111111011111110","0000101111001011110010111100","0000011011110110111101101111","0000011001110110011101100111","0000110100111101001111010011","0000110111001101110011011100","0000011000010110000101100001","0000010011110100111101001111","0000000101110001011100010111","0000010001000100010001000100","0000010011000100110001001100","0000011110010111100101111001","0000100010111000101110001011","0000100011111000111110001111","0000111100111111001111110011","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111100011111000111110001","0000111010001110100011101000","0000011110110111101101111011","0000001101010011010100110101","0000010100010101000101010001","0000001101100011011000110110","0000001100100011001000110010","0000000011110000111100001111","0000001100010011000100110001","0000011111110111111101111111","0000110100101101001011010010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000101111001011110010111100","0000101111101011111010111110","0000110100001101000011010000","0000110101001101010011010100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000110010111100101111001011","0000011110100111101001111010","0000100010111000101110001011","0000011011010110110101101101","0000100000001000000010000000","0000101111001011110010111100","0000111110001111100011111000","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000110010011100100111001001","0000111111111111111111111111","0000111001001110010011100100","0000101011011010110110101101","0001000000000000000000000000","0000100001101000011010000110","0000010011100100111001001110","0000011100100111001001110010","0000100000001000000010000000","0000110101001101010011010100","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110111101101111011011110","0000110001101100011011000110","0000101100001011000010110000","0000101010011010100110101001","0000110000101100001011000010","0000101101001011010010110100","0000110110001101100011011000","0000101010111010101110101011","0000111110111111101111111011","0000110010011100100111001001","0000100001101000011010000110","0000100000011000000110000001","0000000010110000101100001011","0000110011101100111011001110","0000111110101111101011111010","0000110110111101101111011011","0000111001001110010011100100","0000110001001100010011000100","0000110111001101110011011100","0000001100100011001000110010","0000011100100111001001110010","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110",
		"0000111001111110011111100111","0000111110001111100011111000","0000110001111100011111000111","0000000100110001001100010011","0000000011100000111000001110","0000011111100111111001111110","0000100110101001101010011010","0000101010101010101010101010","0000100110101001101010011010","0000101100011011000110110001","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111010011110100111101001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100101111001011110010","0000111101101111011011110110","0000111111011111110111111101","0000110101011101010111010101","0000111101111111011111110111","0000111111001111110011111100","0000111110001111100011111000","0000111000111110001111100011","0000111101111111011111110111","0000111111111111111111111111","0000111101001111010011110100","0000111110001111100011111000","0000111100011111000111110001","0000111111011111110111111101","0000111110101111101011111010","0000011100010111000101110001","0000010111110101111101011111","0000110101111101011111010111","0000110001001100010011000100","0000100110001001100010011000","0000111100011111000111110001","0000111111011111110111111101","0000111110011111100111111001","0000111100011111000111110001","0000111011111110111111101111","0000111111111111111111111111","0000101010111010101110101011","0001000000000000000000000000","0000110001111100011111000111","0000011100000111000001110000","0000100111101001111010011110","0000101010111010101110101011","0000110000011100000111000001","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111110111111101111111011","0000110111101101111011011110","0000101011011010110110101101","0000101001101010011010100110","0000101101101011011010110110","0000110011001100110011001100","0000110010101100101011001010","0000101010001010100010101000","0000100010011000100110001001","0000100001011000010110000101","0000100100001001000010010000","0000100010011000100110001001","0000100011101000111010001110","0000101100101011001010110010","0000110100101101001011010010","0000101011011010110110101101","0000001101110011011100110111","0001000000000000000000000000","0000100010001000100010001000","0000011111000111110001111100","0000011101010111010101110101","0000100010101000101010001010","0000101001111010011110100111","0000101001001010010010100100","0000101111111011111110111111","0000110011001100110011001100","0000110001001100010011000100","0000101010011010100110101001","0000100001001000010010000100","0000100011101000111010001110","0000110001011100010111000101","0000111110101111101011111010","0000110100011101000111010001","0000110100011101000111010001","0000100111101001111010011110","0000011101110111011101110111","0000101100001011000010110000","0000010101010101010101010101","0000010111000101110001011100","0000001101100011011000110110","0000000101000001010000010100","0000001110000011100000111000","0000100101101001011010010110","0000011001100110011001100110","0000100001111000011110000111","0000101111101011111010111110","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111100001111000011110000","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111101111111011111110","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000110111111101111111011111","0000100011011000110110001101","0000011100010111000101110001","0000010110100101101001011010","0000001011010010110100101101","0001000000000000000000000000","0000010010010100100101001001","0000110011111100111111001111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111011101110111011101110","0000101010001010100010101000","0000111100001111000011110000","0000111001011110010111100101","0000111111111111111111111111","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000110001111100011111000111","0000101111011011110110111101","0000100110111001101110011011","0000100111001001110010011100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111100011111000111110001","0000100110011001100110011001","0000010111010101110101011101","0000011001110110011101100111","0000101010001010100010101000","0000100110101001101010011010","0000101111111011111110111111","0000110000111100001111000011","0000111111101111111011111110","0000111111101111111011111110","0000111010111110101111101011","0000110011111100111111001111","0000110010001100100011001000","0000110111111101111111011111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111011001110110011101100","0000110000001100000011000000","0000101110111011101110111011","0000011000000110000001100000","0000100100111001001110010011","0000010111010101110101011101","0000110010111100101111001011","0000100010101000101010001010","0000100001101000011010000110","0000100000001000000010000000","0000011010100110101001101010","0000001010110010101100101011","0000101001001010010010100100","0000110011001100110011001100","0000111101101111011011110110","0000111110111111101111111011","0000111001001110010011100100","0000111001001110010011100100","0000110001111100011111000111","0000001010110010101100101011","0000010101010101010101010101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110111111101111111011","0000101110111011101110111011","0000000010010000100100001001","0000000101000001010000010100","0000011010110110101101101011","0000011001000110010001100100","0000011101110111011101110111","0000100100001001000010010000","0000110010001100100011001000","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111011111110111111101111","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000110001111100011111000111","0000111110001111100011111000","0000111111111111111111111111","0000110100101101001011010010","0000111100011111000111110001","0000111100101111001011110010","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000101101011011010110110101","0000001110010011100100111001","0000101110011011100110111001","0000110010111100101111001011","0000101110001011100010111000","0000110101111101011111010111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000100111101001111010011110","0001000000000000000000000000","0000110101001101010011010100","0000011010110110101101101011","0000011111100111111001111110","0000101010001010100010101000","0000110110011101100111011001","0000111111111111111111111111","0000111100111111001111110011","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111100101111001011110010","0000101011111010111110101111","0000101010011010100110101001","0000100100001001000010010000","0000011101000111010001110100","0000011110000111100001111000","0000100000111000001110000011","0000100001101000011010000110","0000100010111000101110001011","0000101001111010011110100111","0000101110001011100010111000","0000101011001010110010101100","0000011000000110000001100000","0000000100100001001000010010","0000011101100111011001110110","0000101100011011000110110001","0000010011000100110001001100","0000110001001100010011000100","0000101111101011111010111110","0000101011011010110110101101","0000110011101100111011001110","0000101011101010111010101110","0000101111011011110110111101","0000110001011100010111000101","0000101011011010110110101101","0000101110111011101110111011","0000101111001011110010111100","0000100000011000000110000001","0000101101001011010010110100","0000111111111111111111111111","0000110001111100011111000111","0000101110001011100010111000","0000100100011001000110010001","0000100000001000000010000000","0000011000110110001101100011","0000010101110101011101010111","0000001110000011100000111000","0001000000000000000000000000","0000000100110001001100010011","0000101110011011100110111001","0000010000110100001101000011","0000011110110111101101111011","0000100000101000001010000010","0000110000001100000011000000","0000111110101111101011111010","0000111111101111111011111110","0000111101011111010111110101","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111011101110111011101110","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111000111110001111100011","0000010111110101111101011111","0000010111100101111001011110","0000001010110010101100101011","0000001011110010111100101111","0000011100100111001001110010","0000110010011100100111001001","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000101101111011011110110111","0000111100101111001011110010","0000111011011110110111101101","0000111111101111111011111110","0000111111001111110011111100","0000111110001111100011111000","0000111100011111000111110001","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000110001101100011011000110","0000101110001011100010111000","0000100101001001010010010100","0000111100011111000111110001","0000111110111111101111111011","0000111110101111101011111010","0000111100111111001111110011","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000011111010111110101111101","0000010110010101100101011001","0000100001111000011110000111","0000100010111000101110001011","0000100110101001101010011010","0000110000001100000011000000","0000110010101100101011001010","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000101110001011100010111000","0000110010111100101111001011","0000111110011111100111111001","0000111011111110111111101111","0000111110001111100011111000","0000110001001100010011000100","0000111011011110110111101101","0000110000011100000111000001","0000100010101000101010001010","0000001011000010110000101100","0000001100000011000000110000","0000000111010001110100011101","0000011000010110000101100001","0000001011110010111100101111","0000001001010010010100100101","0000000110010001100100011001","0000101010101010101010101010","0000111111111111111111111111","0000111110001111100011111000","0000110011001100110011001100","0000111011001110110011101100","0000111001011110010111100101","0000101011101010111010101110","0000100110001001100010011000","0000010011010100110101001101","0000001111010011110100111101","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111011111110111111101","0000110000111100001111000011","0000000010000000100000001000","0000000010110000101100001011","0000001110110011101100111011","0000001010100010101000101010","0000011011000110110001101100","0000101100111011001110110011","0000111010001110100011101000","0000111101111111011111110111","0000111111101111111011111110","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111110011111100111111001","0000111010101110101011101010","0000101011011010110110101101","0000111010011110100111101001","0000111111111111111111111111","0000101100011011000110110001","0000111101101111011011110110","0000111011111110111111101111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111100001111000011110000","0000111001011110010111100101","0000001110010011100100111001","0000101110011011100110111001","0000111001101110011011100110","0000110000011100000111000001","0000110010011100100111001001","0000111100111111001111110011","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111110001111100011111000","0000100111111001111110011111","0000001000000010000000100000","0000111101001111010011110100","0000011001100110011001100110","0000100110101001101010011010","0000100010001000100010001000","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000111101011111010111110101","0000111101011111010111110101","0000101100011011000110110001","0000101001111010011110100111","0000100011011000110110001101","0000011011000110110001101100","0000010111000101110001011100","0000010011010100110101001101","0000010000110100001101000011","0000011101010111010101110101","0000011110010111100101111001","0000100001011000010110000101","0000100100001001000010010000","0000101000011010000110100001","0000101100101011001010110010","0000100100101001001010010010","0000010100100101001001010010","0000000001110000011100000111","0000101001011010010110100101","0000011011010110110101101101","0000010011010100110101001101","0000101110111011101110111011","0000110000111100001111000011","0000101101001011010010110100","0000110000001100000011000000","0000110111101101111011011110","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000110100001101000011010000","0000101100011011000110110001","0000111011011110110111101101","0000100001111000011110000111","0000110101111101011111010111","0000111011011110110111101101","0000110100101101001011010010","0000101100011011000110110001","0000100011111000111110001111","0000011100100111001001110010","0000011111100111111001111110","0000010101100101011001010110","0001000000000000000000000000","0000000011010000110100001101","0000101000111010001110100011","0000010001110100011101000111","0000011010000110100001101000","0000100100001001000010010000","0000011110110111101101111011","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111110011111100111111001","0000111110011111100111111001","0000111100001111000011110000","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111101101111011011110110","0000111110101111101011111010","0000110000011100000111000001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101100011011000110110001","0000010001000100010001000100","0000000010000000100000001000","0000011110110111101101111011","0000101000001010000010100000","0000110100101101001011010010","0000111101001111010011110100","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111100011111000111110001","0000110011111100111111001111","0000111101001111010011110100","0000111110001111100011111000","0000111111011111110111111101","0000111111011111110111111101","0000111110111111101111111011","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000110011011100110111001101","0000101010011010100110101001","0000110111111101111111011111","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000100000011000000110000001","0000010100000101000001010000","0000100011111000111110001111","0000100001011000010110000101","0000101010001010100010101000","0000110110001101100011011000","0000110010111100101111001011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111010001110100011101000","0000101111011011110110111101","0000100101011001010110010101","0000110110011101100111011001","0000111011001110110011101100","0000110100101101001011010010","0000110011011100110111001101","0000101110101011101010111010","0000101100101011001010110010","0000001110010011100100111001","0001000000000000000000000000","0001000000000000000000000000","0001000000000000000000000000","0000000001110000011100000111","0000011100000111000001110000","0000011010010110100101101001","0000100010101000101010001010","0000101010111010101110101011","0000100101101001011010010110","0000101100011011000110110001","0000101011101010111010101110","0000011000110110001101100011","0000100001111000011110000111","0000011000000110000001100000","0000011100010111000101110001","0000011010000110100001101000","0000110100011101000111010001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111001111110011111100","0000111111001111110011111100","0000110010101100101011001010","0000000001010000010100000101","0000000000110000001100000011","0000000110100001101000011010","0000000110110001101100011011","0000100101011001010110010101","0000111100001111000011110000","0000111111001111110011111100","0000111101111111011111110111","0000111110111111101111111011","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000110010111100101111001011","0000100001111000011110000111","0000110110001101100011011000","0000111011001110110011101100","0000101110001011100010111000","0000110111101101111011011110","0000111100101111001011110010","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000010110110101101101011011","0000101011011010110110101101","0000111000001110000011100000","0000100100111001001110010011","0000111001001110010011100100","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111110011111100111111001","0000111110111111101111111011","0000100111111001111110011111","0000010100010101000101010001","0000111100101111001011110010","0000010000100100001001000010","0000100110011001100110011001","0000101000011010000110100001","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110101111101011111010","0000111111101111111011111110","0000100011111000111110001111","0000100001011000010110000101","0000110000111100001111000011","0000110000001100000011000000","0000011010010110100101101001","0000000001100000011000000110","0000001100010011000100110001","0000000100000001000000010000","0000000001000000010000000100","0000001001010010010100100101","0000010001000100010001000100","0000011010100110101001101010","0000010111100101111001011110","0000001000010010000100100001","0001000000000000000000000000","0001000000000000000000000000","0000000001000000010000000100","0000100000011000000110000001","0000010111110101111101011111","0000011001010110010101100101","0000110010111100101111001011","0000110100111101001111010011","0000111011011110110111101101","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111001111110011111100111","0000111110011111100111111001","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111101101111011011110110","0000110000011100000111000001","0000110111011101110111011101","0000110001011100010111000101","0000111111111111111111111111","0000111101001111010011110100","0000110000101100001011000010","0000100000111000001110000011","0000001110100011101000111010","0000010010010100100101001001","0000010110000101100001011000","0000001111000011110000111100","0001000000000000000000000000","0000010011100100111001001110","0000010110000101100001011000","0000010101000101010001010100","0000101101101011011010110110","0000011011010110110101101101","0000101111101011111010111110","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111101101111011011110110","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000101010111010101110101011","0000110110011101100111011001","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000010010000100100001001000","0001000000000000000000000000","0000100111011001110110011101","0000101100101011001010110010","0000111011111110111111101111","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111101001111010011110100","0000111001111110011111100111","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111000001110000011100000","0000110101011101010111010101","0000110000011100000111000001","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111110011111100111111001","0000111111111111111111111111","0000010101010101010101010101","0000011011100110111001101110","0000100000111000001110000011","0000100001011000010110000101","0000110001011100010111000101","0000111001101110011011100110","0000110101111101011111010111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111001111110011111100","0000111111111111111111111111","0000110001001100010011000100","0000011010100110101001101010","0000100010011000100110001001","0000110101011101010111010101","0000111011111110111111101111","0000101100111011001110110011","0000110100001101000011010000","0000100100101001001010010010","0000011000110110001101100011","0000011011010110110101101101","0000000110010001100100011001","0000000100100001001000010010","0001000000000000000000000000","0001000000000000000000000000","0000000111010001110100011101","0000000010000000100000001000","0000000100010001000100010001","0001000000000000000000000000","0000000010110000101100001011","0000000010000000100000001000","0001000000000000000000000000","0000100000001000000010000000","0000011100000111000001110000","0000010011110100111101001111","0000011001010110010101100101","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000110001001100010011000100","0001000000000000000000000000","0000000011000000110000001100","0000001000010010000100100001","0000001101100011011000110110","0000101111001011110010111100","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000110100001101000011010000","0000100001011000010110000101","0000011000000110000001100000","0000110111101101111011011110","0000101101111011011110110111","0000110101101101011011010110","0000101110011011100110111001","0000111110011111100111111001","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111100101111001011110010","0000011111000111110001111100","0000100111011001110110011101","0000111010001110100011101000","0000011110000111100001111000","0000111100011111000111110001","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111011111110111111101111","0000111111101111111011111110","0000100011101000111010001110","0000011110000111100001111000","0000111010101110101011101010","0000010100010101000101010001","0000011101100111011001110110","0000110000011100000111000001","0000110111101101111011011110","0000111111111111111111111111","0000111110011111100111111001","0000110110101101101011011010","0000011111010111110101111101","0000111001011110010111100101","0000111111001111110011111100","0000101001011010010110100101","0000000011000000110000001100","0000000101000001010000010100","0000010011100100111001001110","0000011011100110111001101110","0000001101010011010100110101","0000010001100100011001000110","0000011010110110101101101011","0000010010000100100001001000","0000010100000101000001010000","0000100010011000100110001001","0000101111101011111010111110","0000111000111110001111100011","0000111101111111011111110111","0000111110011111100111111001","0000110010011100100111001001","0000100001011000010110000101","0000111010111110101111101011","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111110011111100111111001","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100101111001011110010","0000111011011110110111101101","0000101111101011111010111110","0000110001001100010011000100","0000111111011111110111111101","0000111001111110011111100111","0000100011011000110110001101","0000001110000011100000111000","0000010000010100000101000001","0000010010100100101001001010","0000001100110011001100110011","0000000100010001000100010001","0001000000000000000000000000","0000001000100010001000100010","0000011110010111100101111001","0000010010000100100001001000","0000100011001000110010001100","0000100011101000111010001110","0000101001001010010010100100","0000111011111110111111101111","0000111111111111111111111111","0000111100001111000011110000","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100111111001111110011","0000110001011100010111000101","0000100011001000110010001100","0000111101101111011011110110","0000111111011111110111111101","0000111110111111101111111011","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111011011110110111101101","0000100000011000000110000001","0000001000010010000100100001","0000101000101010001010100010","0000101100001011000010110000","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111011001110110011101100","0000111111011111110111111101","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111100101111001011110010","0000111111001111110011111100","0000111110011111100111111001","0000111110011111100111111001","0000111100101111001011110010","0000101011001010110010101100","0000111101101111011011110110","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111100111111001111110011","0000111101101111011011110110","0000111111101111111011111110","0000111001011110010111100101","0000001000100010001000100010","0000101001101010011010100110","0000011011110110111101101111","0000100001011000010110000101","0000110101001101010011010100","0000110111101101111011011110","0000111100001111000011110000","0000111100111111001111110011","0000111110111111101111111011","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000110100101101001011010010","0000100111111001111110011111","0000011111010111110101111101","0000101100111011001110110011","0000110111111101111111011111","0000111011001110110011101100","0000101111001011110010111100","0000101101011011010110110101","0000101000001010000010100000","0000011010100110101001101010","0000011010110110101101101011","0000010110110101101101011011","0000011110010111100101111001","0000101001011010010110100101","0000100111011001110110011101","0000100010001000100010001000","0000011110100111101001111010","0000001111100011111000111110","0000011001010110010101100101","0000100010011000100110001001","0000011011100110111001101110","0000000000010000000100000001","0000000110100001101000011010","0000000110010001100100011001","0000001011100010111000101110","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000000000110000001100000011","0000000111010001110100011101","0000001101010011010100110101","0000010111000101110001011100","0000110010011100100111001001","0000110100111101001111010011","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000110001111100011111000111","0000001100100011001000110010","0000010010000100100001001000","0000111010001110100011101000","0000100001111000011110000111","0000111000011110000111100001","0000101001011010010110100101","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111101111111011111110111","0000111111011111110111111101","0000111111101111111011111110","0000100010111000101110001011","0000011111110111111101111111","0000111111001111110011111100","0000100011101000111010001110","0000111001011110010111100101","0000111110011111100111111001","0000111011111110111111101111","0000111110011111100111111001","0000111011111110111111101111","0000111111001111110011111100","0000011111000111110001111100","0000100010111000101110001011","0000111001111110011111100111","0000100100111001001110010011","0000010101010101010101010101","0000110101001101010011010100","0000111111111111111111111111","0000111101011111010111110101","0000111010011110100111101001","0000101100011011000110110001","0000111101101111011011110110","0000111100001111000011110000","0000110100111101001111010011","0000011001110110011101100111","0000011110110111101101111011","0000011101010111010101110101","0000101000001010000010100000","0000110101111101011111010111","0000101101001011010010110100","0000110011111100111111001111","0000110011011100110111001101","0000110010101100101011001010","0000110100111101001111010011","0000110100001101000011010000","0000101101111011011110110111","0000101100011011000110110001","0000101111111011111110111111","0000110001111100011111000111","0000100100011001000110010001","0000111110101111101011111010","0000111100101111001011110010","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111110011111100111111001","0000111110001111100011111000","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111100111111001111110011","0000111111111111111111111111","0000111110011111100111111001","0000111001111110011111100111","0000100110001001100010011000","0000111110001111100011111000","0000111111111111111111111111","0000110000001100000011000000","0000001000010010000100100001","0000010100110101001101010011","0000010100100101001001010010","0000000001110000011100000111","0000000001100000011000000110","0000001011110010111100101111","0001000000000000000000000000","0000001011010010110100101101","0000010100010101000101010001","0000010010110100101101001011","0000110011011100110111001101","0000101100111011001110110011","0000101000011010000110100001","0000101100001011000010110000","0000110101011101010111010101","0000111100001111000011110000","0000111110001111100011111000","0000111101101111011011110110","0000110100001101000011010000","0000110101011101010111010101","0000101111101011111010111110","0000100001111000011110000111","0000101001101010011010100110","0000110110011101100111011001","0000111001011110010111100101","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000100111111001111110011111","0000001100100011001000110010","0000110100001101000011010000","0000101110001011100010111000","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000110000001100000011000000","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111111101111111011111110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000011110010111100101111001","0000100000111000001110000011","0000101100011011000110110001","0000010100000101000001010000","0000101001111010011110100111","0000110010011100100111001001","0000111000101110001011100010","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000110110001101100011011000","0000010110110101101101011011","0000101101011011010110110101","0000110101101101011011010110","0000111111111111111111111111","0000110100111101001111010011","0000110101111101011111010111","0000101000001010000010100000","0000011101100111011001110110","0000011000000110000001100000","0000011010110110101101101011","0000010111010101110101011101","0000011010100110101001101010","0000100101111001011110010111","0000101011101010111010101110","0000101110101011101010111010","0000110010101100101011001010","0000110010011100100111001001","0000101001111010011110100111","0000010100010101000101010001","0000000110100001101000011010","0000000111000001110000011100","0000000001000000010000000100","0000000111010001110100011101","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101011111010111110101","0000111111111111111111111111","0000101111001011110010111100","0000000010000000100000001000","0000001111010011110100111101","0000010111010101110101011101","0000011111100111111001111110","0000101011011010110110101101","0000110011001100110011001100","0000110100111101001111010011","0000111001111110011111100111","0000111101001111010011110100","0000111110001111100011111000","0000111101111111011111110111","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111110011111100111111001","0000111110111111101111111011","0000101011011010110110101101","0000000001110000011100000111","0000010010110100101101001011","0000110100011101000111010001","0000100000101000001010000010","0000110001111100011111000111","0000101100001011000010110000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000100111001001110010011100","0000010010010100100101001001","0000111010001110100011101000","0000100111111001111110011111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000100001011000010110000101","0000100100101001001010010010","0000110101001101010011010100","0000101100111011001110110011","0000011010000110100001101000","0000110111001101110011011100","0000111101011111010111110101","0000111111111111111111111111","0000110101001101010011010100","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000101100001011000010110000","0000001011110010111100101111","0000011111000111110001111100","0000011111010111110101111101","0000101000001010000010100000","0000111000011110000111100001","0000111000101110001011100010","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111011011110110111101101","0000110011001100110011001100","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111110001111100011111000","0000111110011111100111111001","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111001101110011011100110","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111110101111101011111010","0000110001011100010111000101","0000111010001110100011101000","0000111111111111111111111111","0000111101101111011011110110","0000000111100001111000011110","0000011001110110011101100111","0000010100010101000101010001","0000000110100001101000011010","0000000001110000011100000111","0000000111000001110000011100","0000010011000100110001001100","0000001000110010001100100011","0000000010110000101100001011","0000001011100010111000101110","0000010100110101001101010011","0000010111110101111101011111","0000011111100111111001111110","0000100000011000000110000001","0000011000100110001001100010","0000011000100110001001100010","0000011111000111110001111100","0000100001001000010010000100","0000100010001000100010001000","0000011101100111011001110110","0000100001101000011010000110","0000101101011011010110110101","0000101111011011110110111101","0000111101001111010011110100","0000111100101111001011110010","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111110001111100011111000","0000111011011110110111101101","0000111111111111111111111111","0000100111111001111110011111","0000001111100011111000111110","0000111111101111111011111110","0000110101101101011011010110","0000111001111110011111100111","0000111100111111001111110011","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111000011110000111100001","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000110011111100111111001111","0000010001010100010101000101","0000111010001110100011101000","0000100111111001111110011111","0000011001110110011101100111","0000110011001100110011001100","0000110101111101011111010111","0000111100011111000111110001","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000101100011011000110110001","0000010100000101000001010000","0000011101110111011101110111","0000110111111101111111011111","0000111111111111111111111111","0000111110001111100011111000","0000110111001101110011011100","0000101111011011110110111101","0000101000101010001010100010","0000100000111000001110000011","0000100100001001000010010000","0000101001011010010110100101","0000110001011100010111000101","0000110011011100110111001101","0000111011011110110111101101","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000100111001001110010011100","0000011110010111100101111001","0000000101100001011000010110","0001000000000000000000000000","0000001001000010010000100100","0000110011011100110111001101","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101111111011111110111","0000111101001111010011110100","0000100110101001101010011010","0001000000000000000000000000","0000011000100110001001100010","0000100100111001001110010011","0000100110011001100110011001","0000011111110111111101111111","0000111010101110101011101010","0000110010011100100111001001","0000101100011011000110110001","0000110111111101111111011111","0000111110001111100011111000","0000111001001110010011100100","0000111100001111000011110000","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000100011101000111010001110","0000000001000000010000000100","0000010110010101100101011001","0000101010011010100110101001","0000100101011001010110010101","0000101001111010011110100111","0000110000101100001011000010","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111100001111000011110000","0000111101111111011111110111","0000110000001100000011000000","0000001111100011111000111110","0000111000111110001111100011","0000101001101010011010100110","0000111111111111111111111111","0000111011111110111111101111","0000111111101111111011111110","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000101001001010010010100100","0000101010111010101110101011","0000110101111101011111010111","0000110010011100100111001001","0000011100100111001001110010","0000110101001101010011010100","0000111111101111111011111110","0000110110011101100111011001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000101110011011100110111001","0000000100000001000000010000","0000011110000111100001111000","0000100011011000110110001101","0000110000111100001111000011","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000111100001111000011110000","0000111101011111010111110101","0000111111111111111111111111","0000111101101111011011110110","0000110111101101111011011110","0000111011101110111011101110","0000111010101110101011101010","0000001101010011010100110101","0000010011110100111101001111","0000011100010111000101110001","0001000000000000000000000000","0001000000000000000000000000","0000001100000011000000110000","0000010110000101100001011000","0000001111110011111100111111","0000000001100000011000000110","0001000000000000000000000000","0000001000100010001000100010","0000001001110010011100100111","0000001001100010011000100110","0000001100010011000100110001","0000001100110011001100110011","0000000101110001011100010111","0000001001110010011100100111","0000011010110110101101101011","0000100011111000111110001111","0000101001001010010010100100","0000101111001011110010111100","0000110110101101101011011010","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111101101111011011110110","0000111111011111110111111101","0000111110011111100111111001","0000111011001110110011101100","0000111011001110110011101100","0000101011011010110110101101","0000011000110110001101100011","0000111110011111100111111001","0000111101011111010111110101","0000110000111100001111000011","0000111011101110111011101110","0000111111111111111111111111","0000111100011111000111110001","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000110101011101010111010101","0000011111110111111101111111","0000011111100111111001111110","0000110010001100100011001000","0000100111111001111110011111","0000101100011011000110110001","0000110011001100110011001100","0000111111101111111011111110","0000111100001111000011110000","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111110101111101011111010","0000111101101111011011110110","0000111110001111100011111000","0000111111101111111011111110","0000111111101111111011111110","0000010111010101110101011101","0000010110110101101101011011","0000100100011001000110010001","0000111110111111101111111011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111001001110010011100100","0000111011001110110011101100","0000110100001101000011010000","0000110011011100110111001101","0000110110111101101111011011","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111011011110110111101101","0000111111011111110111111101","0000111100101111001011110010","0000010111110101111101011111","0000001001000010010000100100","0000000000010000000100000001","0000000110000001100000011000","0000101101111011011110110111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110011111100111111001","0000001110100011101000111010","0001000000000000000000000000","0000101010101010101010101010","0000111001011110010111100101","0000101100001011000010110000","0000100101101001011010010110","0000101010101010101010101010","0000111011001110110011101100","0000111101101111011011110110","0000100110111001101110011011","0000101101111011011110110111","0000111110111111101111111011","0000111010001110100011101000","0000101111101011111010111110","0000111000011110000111100001","0000111011001110110011101100","0000110011111100111111001111","0000001110010011100100111001","0000000010100000101000001010","0000100000111000001110000011","0000100101011001010110010101","0000010111000101110001011100","0000100010011000100110001001","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000110010001100100011001000","0000000110100001101000011010","0000110111111101111111011111","0000101101111011011110110111","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000101110101011101010111010","0000110011011100110111001101","0000111011101110111011101110","0000111101111111011111110111","0000100010101000101010001010","0000111001101110011011100110","0000111111111111111111111111","0000111100101111001011110010","0000111101001111010011110100","0000111110111111101111111011","0000111100111111001111110011","0000011110110111101101111011","0000001100100011001000110010","0000100110011001100110011001","0000110110101101101011011010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111110001111100011111000","0000111101101111011011110110","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111110001111100011111000","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111100001111000011110000","0000111110111111101111111011","0000111110001111100011111000","0000111010011110100111101001","0000111111111111111111111111","0000111100101111001011110010","0000001010100010101000101010","0000001001100010011000100110","0000010001000100010001000100","0000000000010000000100000001","0001000000000000000000000000","0000010011110100111101001111","0000001100100011001000110010","0001000000000000000000000000","0000001011110010111100101111","0000010010110100101101001011","0000011011010110110101101101","0000100001011000010110000101","0000100000001000000010000000","0000011100000111000001110000","0000011101000111010001110100","0000100011101000111010001110","0000011110000111100001111000","0000010011100100111001001110","0000100011001000110010001100","0000111011001110110011101100","0000111111111111111111111111","0000111100101111001011110010","0000111100101111001011110010","0000111111111111111111111111","0000111011001110110011101100","0000111110101111101011111010","0000111111101111111011111110","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000110001001100010011000100","0000110001001100010011000100","0000010001110100011101000111","0000111010001110100011101000","0000111000001110000011100000","0000110011001100110011001100","0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111111101111111011111110","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111110001111100011111000","0000111101111111011111110111","0000111011111110111111101111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111001111110011111100111","0000101011011010110110101101","0000010111000101110001011100","0000000110000001100000011000","0000101011101010111010101110","0000101111001011110010111100","0000111001111110011111100111","0000101010011010100110101001","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000011111110111111101111111","0001000000000000000000000000","0000100111001001110010011100","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111010111110101111101011","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000101100001011000010110000","0000000101010001010100010101","0000001111000011110000111100","0000000010100000101000001010","0000101011111010111110101111","0000111111111111111111111111","0000111110101111101011111010",
		"0000111101011111010111110101","0000111010111110101111101011","0000001000000010000000100000","0000000011110000111100001111","0000110000111100001111000011","0000111100111111001111110011","0000110110001101100011011000","0000101110101011101010111010","0000100000001000000010000000","0000101010001010100010101000","0000111010001110100011101000","0000110111001101110011011100","0000101000001010000010100000","0000100000001000000010000000","0000101111001011110010111100","0000111010001110100011101000","0000100001101000011010000110","0000011100000111000001110000","0000101010001010100010101000","0000010001100100011001000110","0000000111110001111100011111","0000011010100110101001101010","0000011101110111011101110111","0000010100010101000101010001","0000100111001001110010011100","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000110100111101001111010011","0000000011110000111100001111","0000111000111110001111100011","0000101110111011101110111011","0000111111011111110111111101","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111110011111100111111001","0000111010111110101111101011","0000100111011001110110011101","0000110110101101101011011010","0000111100101111001011110010","0000111011011110110111101101","0000101010101010101010101010","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111010111110101111101011","0000110010011100100111001001","0000101000001010000010100000","0000011011100110111001101110","0000110001101100011011000110","0000111100111111001111110011","0000111111101111111011111110","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111100001111000011110000","0000111011011110110111101101","0000111101011111010111110101","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111111011111110111111101","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111011011110110111101101","0000111100011111000111110001","0000110110001101100011011000","0000000100000001000000010000","0000001101100011011000110110","0000010100010101000101010001","0000000001010000010100000101","0000000001010000010100000101","0000000101000001010000010100","0000001001100010011000100110","0000010000110100001101000011","0000010101010101010101010101","0000001011010010110100101101","0000010001010100010101000101","0000010101000101010001010100","0000011100000111000001110000","0000011100010111000101110001","0000100010101000101010001010","0000100010111000101110001011","0000100100101001001010010010","0000100001001000010010000100","0000101011101010111010101110","0000101110001011100010111000","0000110111011101110111011101","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111001001110010011100100","0000110001001100010011000100","0000110000111100001111000011","0000001011110010111100101111","0000101010101010101010101010","0000101101001011010010110100","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111011101110111011101110","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111100101111001011110010","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111001111110011111100111","0000111111111111111111111111","0000111001111110011111100111","0000111101001111010011110100","0000111111111111111111111111","0000111010101110101011101010","0000111100111111001111110011","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110100001101000011010000","0000010001100100011001000110","0000010110000101100001011000","0000000011010000110100001101","0000011010110110101101101011","0000111101111111011111110111","0000110000111100001111000011","0000101101101011011010110110","0000110001011100010111000101","0000111110101111101011111010","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000110001011100010111000101","0000000001100000011000000110","0000010001110100011101000111","0000110100001101000011010000","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000110101001101010011010100","0000001100110011001100110011","0000010100000101000001010000","0001000000000000000000000000","0000100001011000010110000101","0000111111111111111111111111","0000111110111111101111111011",
		"0000111011111110111111101111","0000110110111101101111011011","0000000001100000011000000110","0000001010110010101100101011","0000111000011110000111100001","0000111111111111111111111111","0000111111101111111011111110","0000111000011110000111100001","0000101111111011111110111111","0000011110110111101101111011","0000011111110111111101111111","0000110101001101010011010100","0000101111101011111010111110","0000100101001001010010010100","0000000111000001110000011100","0000001100110011001100110011","0000011010110110101101101011","0000100000001000000010000000","0000010110010101100101011001","0000000010110000101100001011","0000010010010100100101001001","0000011011110110111101101111","0000010111100101111001011110","0000010011010100110101001101","0000101101011011010110110101","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111110111111101111111011","0000111110001111100011111000","0000111111101111111011111110","0000110111011101110111011101","0000000100000001000000010000","0000110111001101110011011100","0000110011001100110011001100","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111111111111111111111111","0000111100001111000011110000","0000111001011110010111100101","0000100101001001010010010100","0000111011101110111011101110","0000111111101111111011111110","0000110111111101111111011111","0000110011101100111011001110","0000111000111110001111100011","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100001101000011010000","0000110010111100101111001011","0000101101011011010110110101","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111110111111101111111011","0000111110011111100111111001","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100011111000111110001","0000111111111111111111111111","0000111101101111011011110110","0000110111001101110011011100","0000111100101111001011110010","0000111011011110110111101101","0000111111111111111111111111","0000111010101110101011101010","0000111111001111110011111100","0000111111111111111111111111","0000101111101011111010111110","0000000100110001001100010011","0000001110010011100100111001","0000001011000010110000101100","0000000101100001011000010110","0001000000000000000000000000","0000000001100000011000000110","0000011100110111001101110011","0000011110100111101001111010","0000010011110100111101001111","0000010000110100001101000011","0000010010100100101001001010","0000100000101000001010000010","0000011111100111111001111110","0000011011100110111001101110","0000011010110110101101101011","0000101010101010101010101010","0000100010111000101110001011","0000010011010100110101001101","0000011111010111110101111101","0000110011011100110111001101","0000111111011111110111111101","0000111011011110110111101101","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000110110001101100011011000","0000110000101100001011000010","0000101001011010010110100101","0000000111000001110000011100","0000100111111001111110011111","0000101110111011101110111011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000110111111101111111011111","0000111000001110000011100000","0000101100111011001110110011","0000101011101010111010101110","0000101001001010010010100100","0000101001011010010110100101","0000100111101001111010011110","0000100111111001111110011111","0000101000101010001010100010","0000100100111001001110010011","0000100011001000110010001100","0000100111011001110110011101","0000101011001010110010101100","0000100000001000000010000000","0000011000010110000101100001","0000010110010101100101011001","0000000100010001000100010001","0000001100010011000100110001","0000011001100110011001100110","0000111110001111100011111000","0000110111011101110111011101","0000101101001011010010110100","0000101001011010010110100101","0000111010001110100011101000","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000000110100001101000011010","0000000001010000010100000101","0000100011011000110110001101","0000111101001111010011110100","0000111110001111100011111000","0000111100101111001011110010","0000111111011111110111111101","0000111100101111001011110010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111001101110011011100110","0000111001111110011111100111","0000111111101111111011111110","0000111111111111111111111111","0000111100101111001011110010","0000111000111110001111100011","0000100100011001000110010001","0000100110011001100110011001","0000010111010101110101011101","0001000000000000000000000000","0000010001000100010001000100","0000111111111111111111111111","0000111111001111110011111100",
		"0000111110011111100111111001","0000110011001100110011001100","0001000000000000000000000000","0000010001100100011001000110","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110001101100011011000110","0000100100011001000110010001","0000011011100110111001101110","0000011100010111000101110001","0000100010101000101010001010","0000101001011010010110100101","0000110011101100111011001110","0000100001001000010010000100","0000001010010010100100101001","0000011011100110111001101110","0000011110000111100001111000","0000010011000100110001001100","0000011000100110001001100010","0000011011000110110001101100","0000010101010101010101010101","0000010011110100111101001111","0000110001101100011011000110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111010011110100111101001","0000001000010010000100100001","0000110010101100101011001010","0000111001001110010011100100","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111000101110001011100010","0000111001001110010011100100","0000101001001010010010100100","0000111111101111111011111110","0000111111111111111111111111","0000110111011101110111011101","0000110001101100011011000110","0000111001011110010111100101","0000111111011111110111111101","0000111111111111111111111111","0000111101011111010111110101","0000110111001101110011011100","0000110010111100101111001011","0000110000101100001011000010","0000110110011101100111011001","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111100001111000011110000","0000111100011111000111110001","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000110111011101110111011101","0000110010101100101011001010","0000101100011011000110110001","0000100011001000110010001100","0000100000001000000010000000","0000100010011000100110001001","0000100101011001010110010101","0000101001101010011010100110","0000101011101010111010101110","0000101010011010100110101001","0000101101011011010110110101","0000110100011101000111010001","0000111111111111111111111111","0000110111101101111011011110","0000110000001100000011000000","0000001110010011100100111001","0000010000000100000001000000","0000001001110010011100100111","0000001011100010111000101110","0000000011100000111000001110","0000000001110000011100000111","0000010010010100100101001001","0000010101000101010001010100","0000001111010011110100111101","0000011111010111110101111101","0000100010001000100010001000","0000100000101000001010000010","0000100110111001101110011011","0000110010101100101011001010","0000110000001100000011000000","0000110100101101001011010010","0000101111111011111110111111","0000110011101100111011001110","0000110001001100010011000100","0000101100101011001010110010","0000101011011010110110101101","0000110101011101010111010101","0000111111111111111111111111","0000111100011111000111110001","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000110110111101101111011011","0000101010101010101010101010","0000100110101001101010011010","0000001011110010111100101111","0000100111001001110010011100","0000110010111100101111001011","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111111011111110111111101","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111011101110111011101110","0000011001110110011101100111","0000110010011100100111001001","0000110011001100110011001100","0000110111101101111011011110","0000110111101101111011011110","0000100001011000010110000101","0000010001100100011001000110","0000001110000011100000111000","0000010001010100010101000101","0000010001000100010001000100","0000011001110110011101100111","0000100101011001010110010101","0000100101111001011110010111","0000011000010110000101100001","0000010001100100011001000110","0001000000000000000000000000","0000010001000100010001000100","0000010100010101000101010001","0000010100110101001101010011","0000111001011110010111100101","0000111001101110011011100110","0000101011111010111110101111","0000101010001010100010101000","0000101111111011111110111111","0000111110101111101011111010","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000010111110101111101011111","0000001010000010100000101000","0000011100110111001101110011","0000110011001100110011001100","0000111001001110010011100100","0000111110111111101111111011","0000111111101111111011111110","0000111101111111011111110111","0000111100001111000011110000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111001101110011011100110","0000101110001011100010111000","0000100110101001101010011010","0000111111111111111111111111","0000101110111011101110111011","0000101000001010000010100000","0001000000000000000000000000","0000001000000010000000100000","0000111011101110111011101110","0000111111011111110111111101",
		"0000111111111111111111111111","0000101110111011101110111011","0001000000000000000000000000","0000010110110101101101011011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000110111001101110011011100","0000101010101010101010101010","0000100011111000111110001111","0000100001101000011010000110","0000011100110111001101110011","0000010000110100001101000011","0000100001001000010010000100","0000100010101000101010001010","0000010010000100100001001000","0000001010000010100000101000","0000011101100111011001110110","0000000011000000110000001100","0000100101011001010110010101","0000010111110101111101011111","0000010000100100001001000010","0000110000111100001111000011","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000001101010011010100110101","0000101110011011100110111001","0000111011011110110111101101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000101101011011010110110101","0000110101101101011011010110","0000101001001010010010100100","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111001101110011011100110","0000111000001110000011100000","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111000011110000111100001","0000111100101111001011110010","0000101010011010100110101001","0000111001001110010011100100","0000111111111111111111111111","0000111100111111001111110011","0000111100011111000111110001","0000111111011111110111111101","0000111111001111110011111100","0000111111011111110111111101","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000101111101011111010111110","0000100010111000101110001011","0000011100000111000001110000","0000011110000111100001111000","0000100110011001100110011001","0000101101101011011010110110","0000101100011011000110110001","0000101010101010101010101010","0000101000101010001010100010","0000101010001010100010101000","0000101101001011010010110100","0000101110011011100110111001","0000101010001010100010101000","0000100001111000011110000111","0000100001001000010010000100","0000100010101000101010001010","0000100111101001111010011110","0000100000111000001110000011","0000011011100110111001101110","0000010001010100010101000101","0000001011010010110100101101","0000010000100100001001000010","0000010000010100000101000001","0001000000000000000000000000","0000000000110000001100000011","0000010100000101000001010000","0000010101100101011001010110","0000010100000101000001010000","0000100110001001100010011000","0000011100000111000001110000","0000101011001010110010101100","0000101011001010110010101100","0000101110111011101110111011","0000111111111111111111111111","0000111100101111001011110010","0000111001011110010111100101","0000110101001101010011010100","0000111110101111101011111010","0000110011011100110111001101","0000110101101101011011010110","0000110000111100001111000011","0000110110101101101011011010","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111111101111111011111110","0000111101111111011111110111","0000111110111111101111111011","0000110110101101101011011010","0000011110000111100001111000","0000100110001001100010011000","0000010001010100010101000101","0000010101010101010101010101","0000110101011101010111010101","0000111101101111011011110110","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110111111101111111011111","0000100010001000100010001000","0000111110011111100111111001","0000111101001111010011110100","0000111101011111010111110101","0000100001111000011110000111","0000000011000000110000001100","0000000010010000100100001001","0000000000110000001100000011","0000001010000010100000101000","0000001111100011111000111110","0000000111110001111100011111","0000000111010001110100011101","0000010001110100011101000111","0000011000010110000101100001","0000011100110111001101110011","0000100000101000001010000010","0000010111010101110101011101","0000011011110110111101101111","0000001101000011010000110100","0000110110111101101111011011","0000101010011010100110101001","0000110010011100100111001001","0000101110101011101010111010","0000101101011011010110110101","0000111000111110001111100011","0000111110101111101011111010","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111011011110110111101101","0000010001100100011001000110","0000000110000001100000011000","0000100101011001010110010101","0000111000011110000111100001","0000101011101010111010101110","0000101100101011001010110010","0000110100011101000111010001","0000110111001101110011011100","0000111000011110000111100001","0000110111011101110111011101","0000110110111101101111011011","0000110110001101100011011000","0000110010101100101011001010","0000101101111011011110110111","0000100011001000110010001100","0000110110111101101111011011","0000111111011111110111111101","0000111011101110111011101110","0000110011111100111111001111","0000101010101010101010101010","0000010001000100010001000100","0000010000010100000101000001","0000110000101100001011000010","0000111111111111111111111111",
		"0000111111111111111111111111","0000101101001011010010110100","0001000000000000000000000000","0000011011010110110101101101","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000110100101101001011010010","0000100000001000000010000000","0000011000110110001101100011","0000001001010010010100100101","0000011010010110100101101001","0000011000110110001101100011","0000011110100111101001111010","0000100001101000011010000110","0000001011100010111000101110","0000010110100101101001011010","0000001010100010101000101010","0000010011100100111001001110","0000010110000101100001011000","0000010111110101111101011111","0000101011011010110110101101","0000111101011111010111110101","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000010011000100110001001100","0000100111101001111010011110","0000111010001110100011101000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000110101001101010011010100","0000100000101000001010000010","0000101101001011010010110100","0000100111001001110010011100","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000110101001101010011010100","0000110010001100100011001000","0000111100101111001011110010","0000111111111111111111111111","0000111101111111011111110111","0000101101101011011010110110","0000111100111111001111110011","0000101111011011110110111101","0000111011001110110011101100","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000110010011100100111001001","0000110101101101011011010110","0000111010001110100011101000","0000111101001111010011110100","0000111101011111010111110101","0000111010111110101111101011","0000110111111101111111011111","0000110101111101011111010111","0000101001101010011010100110","0000100010111000101110001011","0000001000110010001100100011","0001000000000000000000000000","0000010000000100000001000000","0000011001010110010101100101","0000011000010110000101100001","0000011001000110010001100100","0000011010100110101001101010","0000010100100101001001010010","0000100000111000001110000011","0000100100001001000010010000","0000011100000111000001110000","0000010001110100011101000111","0000011110100111101001111010","0000011000100110001001100010","0000001100000011000000110000","0000000001000000010000000100","0000000100000001000000010000","0000000110100001101000011010","0000001011110010111100101111","0000010101000101010001010100","0000100111101001111010011110","0000110010001100100011001000","0000110111011101110111011101","0000110110101101101011011010","0000111001111110011111100111","0000110110111101101111011011","0000111111111111111111111111","0000111110111111101111111011","0000111011001110110011101100","0000101111011011110110111101","0000111011101110111011101110","0000110010111100101111001011","0000110110101101101011011010","0000111010111110101111101011","0000111101011111010111110101","0000111010101110101011101010","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111100001111000011110000","0000111111101111111011111110","0000111010111110101111101011","0000010011100100111001001110","0000011001010110010101100101","0000010000010100000101000001","0000001000000010000000100000","0000110001001100010011000100","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000110000011100000111000001","0000100011011000110110001101","0000111101011111010111110101","0000111110101111101011111010","0000110110101101101011011010","0000001110010011100100111001","0000000011000000110000001100","0000100101011001010110010101","0000101110101011101010111010","0000101111011011110110111101","0000101011101010111010101110","0000101101001011010010110100","0000101101101011011010110110","0000011001110110011101100111","0000000011110000111100001111","0000000000100000001000000010","0000010001010100010101000101","0000100000001000000010000000","0000100001001000010010000100","0000010111000101110001011100","0000100011101000111010001110","0000110000001100000011000000","0000101101111011011110110111","0000110001011100010111000101","0000100110001001100010011000","0000110010001100100011001000","0000111111111111111111111111","0000111110101111101011111010","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111000011110000111100001","0000011101000111010001110100","0000001011100010111000101110","0000100010111000101110001011","0000110001011100010111000101","0000101011011010110110101101","0000101010011010100110101001","0000100101011001010110010101","0000100011011000110110001101","0000100100001001000010010000","0000100111001001110010011100","0000101000001010000010100000","0000100111111001111110011111","0000101011001010110010101100","0000110000001100000011000000","0000111001001110010011100100","0000101110111011101110111011","0000111000001110000011100000","0000111100001111000011110000","0000111000001110000011100000","0000101011101010111010101110","0000011110110111101101111011","0000011000010110000101100001","0000100001011000010110000101","0000111111111111111111111111",
		"0000111111111111111111111111","0000110000011100000111000001","0001000000000000000000000000","0000100000011000000110000001","0000111100011111000111110001","0000111001111110011111100111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110001111100011111000","0000111010101110101011101010","0000110000111100001111000011","0000100001001000010010000100","0000011111000111110001111100","0000011010010110100101101001","0000100111101001111010011110","0000011001110110011101100111","0000000100100001001000010010","0000011010110110101101101011","0000000001110000011100000111","0000011001110110011101100111","0000101100101011001010110010","0000100100001001000010010000","0000111000101110001011100010","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111110101111101011111010","0000011101000111010001110100","0000011010110110101101101011","0000111011001110110011101100","0000110110011101100111011001","0000111111011111110111111101","0000111111111111111111111111","0000101111011011110110111101","0000011110010111100101111001","0000100011101000111010001110","0000101110111011101110111011","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110011101100111011001110","0000111010111110101111101011","0000110001001100010011000100","0000110101111101011111010111","0000111111001111110011111100","0000111110101111101011111010","0000111110001111100011111000","0000111101101111011011110110","0000111011011110110111101101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111101101111011011110110","0000111100111111001111110011","0000111010001110100011101000","0000110100111101001111010011","0000110000111100001111000011","0000110000101100001011000010","0000100111111001111110011111","0000001010000010100000101000","0001000000000000000000000000","0000001100110011001100110011","0000001011110010111100101111","0000000011010000110100001101","0000000001010000010100000101","0000010010110100101101001011","0000011110000111100001111000","0000010100110101001101010011","0000100111101001111010011110","0000101011111010111110101111","0000100110011001100110011001","0000100100011001000110010001","0000011010000110100001101000","0000000110100001101000011010","0000000011000000110000001100","0000000001010000010100000101","0000001111010011110100111101","0000001110010011100100111001","0000100111011001110110011101","0000101100111011001110110011","0000101111011011110110111101","0000110001001100010011000100","0000111001101110011011100110","0000111100101111001011110010","0000111110111111101111111011","0000111011111110111111101111","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000110101101101011011010110","0000111111111111111111111111","0000111101011111010111110101","0000110001011100010111000101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111011001110110011101100","0000001111110011111100111111","0000001111110011111100111111","0000011000000110000001100000","0000001110100011101000111010","0000100001011000010110000101","0000101100011011000110110001","0000111000111110001111100011","0000111100011111000111110001","0000111110101111101011111010","0000111001111110011111100111","0000101110011011100110111001","0000100111011001110110011101","0000101000101010001010100010","0000111111111111111111111111","0000110001111100011111000111","0000100111111001111110011111","0001000000000000000000000000","0000011000100110001001100010","0000111001111110011111100111","0000111100001111000011110000","0000111001001110010011100100","0000101101111011011110110111","0000100111001001110010011100","0000100100111001001110010011","0000011100010111000101110001","0000010000000100000001000000","0000001000110010001100100011","0000000111010001110100011101","0000000110110001101100011011","0000001010010010100100101001","0000001101100011011000110110","0000011101100111011001110110","0000101101101011011010110110","0000101100001011000010110000","0000100110001001100010011000","0000100111111001111110011111","0000100100101001001010010010","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110010101100101011001010","0000101010001010100010101000","0000100001111000011110000111","0000001110000011100000111000","0000100111001001110010011100","0000101000011010000110100001","0000100101011001010110010101","0000011101100111011001110110","0000011111010111110101111101","0000011000100110001001100010","0000001100000011000000110000","0000000101000001010000010100","0000001111100011111000111110","0000100010011000100110001001","0000101010011010100110101001","0000100111011001110110011101","0000110100111101001111010011","0000111001011110010111100101","0000111111111111111111111111","0000111101101111011011110110","0000111011101110111011101110","0000101011101010111010101110","0000011100000111000001110000","0000100101101001011010010110","0000010010010100100101001001","0000111111111111111111111111",
		"0000111111111111111111111111","0000110101101101011011010110","0001000000000000000000000000","0000100100001001000010010000","0000111100001111000011110000","0000110101001101010011010100","0000111111111111111111111111","0000111010111110101111101011","0000111110011111100111111001","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000110111001101110011011100","0000101111001011110010111100","0000011010110110101101101011","0000011001010110010101100101","0000011010110110101101101011","0000000000110000001100000011","0000001111000011110000111100","0000001100100011001000110010","0000110100011101000111010001","0000011110110111101101111011","0000110101101101011011010110","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111100011111000111110001","0000111000101110001011100010","0000100110101001101010011010","0000001110100011101000111010","0000111101111111011111110111","0000101111101011111010111110","0000111111001111110011111100","0000111100101111001011110010","0000101010011010100110101001","0000100011111000111110001111","0000011101100111011001110110","0000111011011110110111101101","0000111100001111000011110000","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111010101110101011101010","0000111111001111110011111100","0000111101111111011111110111","0000111101011111010111110101","0000110111101101111011011110","0000111010001110100011101000","0000111001101110011011100110","0000101010101010101010101010","0000110110111101101111011011","0000111001001110010011100100","0000111000001110000011100000","0000110101001101010011010100","0000110010111100101111001011","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000110111011101110111011101","0000110100001101000011010000","0000110010101100101011001010","0000111000011110000111100001","0000110111001101110011011100","0000101111001011110010111100","0000101110011011100110111001","0000101001001010010010100100","0000010111100101111001011110","0000001010100010101000101010","0000000001110000011100000111","0001000000000000000000000000","0000001011110010111100101111","0000010111000101110001011100","0000011010000110100001101000","0000101011011010110110101101","0000101111011011110110111101","0000101101101011011010110110","0000100110111001101110011011","0001000000000000000000000000","0000100000001000000010000000","0001000000000000000000000000","0000010001110100011101000111","0000010100100101001001010010","0000110100111101001111010011","0000100110001001100010011000","0000101100001011000010110000","0000110100111101001111010011","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000110111011101110111011101","0000111111001111110011111100","0000111011011110110111101101","0000111010111110101111101011","0000111100101111001011110010","0000111111011111110111111101","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110010111100101111001011","0000001111110011111100111111","0000010101110101011101010111","0000101001101010011010100110","0000010111110101111101011111","0000011001000110010001100100","0000100001001000010010000100","0000100100111001001110010011","0000100110001001100010011000","0000100011011000110110001101","0000100000011000000110000001","0000011010010110100101101001","0000101001111010011110100111","0000110001001100010011000100","0000100100011001000110010001","0000010001100100011001000110","0001000000000000000000000000","0000101111001011110010111100","0000111111101111111011111110","0000111110011111100111111001","0000111100011111000111110001","0000111001001110010011100100","0000111010101110101011101010","0000101111101011111010111110","0000101000111010001110100011","0000100111001001110010011100","0000010101110101011101010111","0000001011000010110000101100","0000010111010101110101011101","0000010101010101010101010101","0001000000000000000000000000","0000000101010001010100010101","0000010001000100010001000100","0000101101001011010010110100","0000011000100110001001100010","0000101100011011000110110001","0000011010010110100101101001","0000111010001110100011101000","0000111111111111111111111111","0000110111001101110011011100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000011111010111110101111101","0000100101011001010110010101","0000101011001010110010101100","0000010111000101110001011100","0000111100101111001011110010","0000100100101001001010010010","0000010110000101100001011000","0000010110110101101101011011","0000000001100000011000000110","0000000001010000010100000101","0000000010110000101100001011","0000001000110010001100100011","0000010110000101100001011000","0000100111101001111010011110","0000110111011101110111011101","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111111011111110111111101","0000111101111111011111110111","0000111111011111110111111101","0000110010101100101011001010","0000100001101000011010000110","0000101101001011010010110100","0000001000110010001100100011","0000111111111111111111111111",
		"0000111110111111101111111011","0000111100111111001111110011","0000001000000010000000100000","0000011111100111111001111110","0000111011011110110111101101","0000110000011100000111000001","0000111110111111101111111011","0000110111101101111011011110","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000110111001101110011011100","0000110111011101110111011101","0000111111111111111111111111","0000111110011111100111111001","0000111100001111000011110000","0000111010111110101111101011","0000100110011001100110011001","0000101101111011011110110111","0000010011000100110001001100","0000001111100011111000111110","0000010100010101000101010001","0000101000011010000110100001","0000110000111100001111000011","0000100110001001100010011000","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111000111110001111100011","0000111111101111111011111110","0000111111101111111011111110","0000111110001111100011111000","0000111001111110011111100111","0000100011011000110110001101","0000000101100001011000010110","0000110111001101110011011100","0000100010101000101010001010","0000111111111111111111111111","0000111110001111100011111000","0000100010111000101110001011","0000101000111010001110100011","0000011011110110111101101111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111010101110101011101010","0000111110101111101011111010","0000101100001011000010110000","0000100000001000000010000000","0000101111011011110110111101","0000110101001101010011010100","0000100000111000001110000011","0000101000111010001110100011","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111100111111001111110011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111001001110010011100100","0000110000011100000111000001","0000101000111010001110100011","0000101001001010010010100100","0000101011111010111110101111","0000100111101001111010011110","0000011111010111110101111101","0000000110110001101100011011","0000001001110010011100100111","0000101000001010000010100000","0000011100000111000001110000","0000010011010100110101001101","0000011010010110100101101001","0000110011101100111011001110","0000110000111100001111000011","0000000001110000011100000111","0000100111101001111010011110","0001000000000000000000000000","0000001001110010011100100111","0000011111000111110001111100","0000110100001101000011010000","0000100001011000010110000101","0000101000011010000110100001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111011111110111111101","0000111100111111001111110011","0000111101001111010011110100","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111110001111100011111000","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111100011111000111110001","0000111110001111100011111000","0000110010101100101011001010","0000011010010110100101101001","0000100001011000010110000101","0000110011111100111111001111","0000100011001000110010001100","0000010001010100010101000101","0000010101110101011101010111","0000010010010100100101001001","0000001011100010111000101110","0000010011010100110101001101","0000010011000100110001001100","0000011111110111111101111111","0000010011110100111101001111","0001000000000000000000000000","0000000011100000111000001110","0000011011100110111001101110","0000110111001101110011011100","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111001101110011011100110","0000101101111011011110110111","0000010100000101000001010000","0001000000000000000000000000","0000000001000000010000000100","0000000110100001101000011010","0000010001100100011001000110","0000100000101000001010000010","0000011100110111001101110011","0000110000101100001011000010","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111010011110100111101001","0000111111111111111111111111","0000111101011111010111110101","0000111101101111011011110110","0000111111111111111111111111","0000101010101010101010101010","0000100000101000001010000010","0000101100001011000010110000","0000110010101100101011001010","0000001101110011011100110111","0000100001111000011110000111","0000000010100000101000001010","0001000000000000000000000000","0000011000100110001001100010","0000101101011011010110110101","0000110000011100000111000001","0000110101001101010011010100","0000111001111110011111100111","0000111101011111010111110101","0000111110111111101111111011","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000110111001101110011011100","0000100010101000101010001010","0000111000101110001011100010","0000001000000010000000100000","0000111001111110011111100111",
		"0000111110101111101011111010","0000111101001111010011110100","0000000110110001101100011011","0000011111010111110101111101","0000110000011100000111000001","0000101100111011001110110011","0000111101101111011011110110","0000110011001100110011001100","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000101010001010100010101000","0000111010111110101111101011","0000111110001111100011111000","0000111111101111111011111110","0000111011101110111011101110","0000110011111100111111001111","0000111111101111111011111110","0000100110101001101010011010","0000100011111000111110001111","0000000111000001110000011100","0000011100010111000101110001","0000100001001000010010000100","0000111010111110101111101011","0000011010010110100101101001","0000110101111101011111010111","0000111111111111111111111111","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111101011111010111110101","0000111101101111011011110110","0000111111101111111011111110","0000111101111111011111110111","0000101110111011101110111011","0000000000110000001100000011","0000100111101001111010011110","0000111000011110000111100001","0000101010101010101010101010","0000111111111111111111111111","0000100011001000110010001100","0000100000001000000010000000","0000011110010111100101111001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111011001110110011101100","0000111111111111111111111111","0000111100111111001111110011","0000111110001111100011111000","0000111111101111111011111110","0000111101101111011011110110","0000101111001011110010111100","0000100111101001111010011110","0000011111110111111101111111","0000101100001011000010110000","0000101001101010011010100110","0000101000001010000010100000","0000111101101111011011110110","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110001111100011111000","0000110111111101111111011111","0000101011101010111010101110","0000100010101000101010001010","0000100000101000001010000010","0000100000001000000010000000","0000011110000111100001111000","0000100110001001100010011000","0000010110110101101101011011","0000000000100000001000000010","0000101010001010100010101000","0000100110101001101010011010","0000010010100100101001001010","0000010111110101111101011111","0000110011011100110111001101","0001000000000000000000000000","0000100101101001011010010110","0000000001000000010000000100","0000000011000000110000001100","0000100000011000000110000001","0000011101100111011001110110","0000011011010110110101101101","0000101110011011100110111001","0000111110101111101011111010","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111010101110101011101010","0000111110111111101111111011","0000111011101110111011101110","0000111110011111100111111001","0000111111101111111011111110","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000110110111101101111011011","0000110001111100011111000111","0000101110111011101110111011","0000100000001000000010000000","0000010101010101010101010101","0000011000010110000101100001","0000101000001010000010100000","0000011100110111001101110011","0000011100010111000101110001","0000101000001010000010100000","0000011100010111000101110001","0000100010001000100010001000","0000010110000101100001011000","0000010110100101101001011010","0001000000000000000000000000","0000000010100000101000001010","0000001011110010111100101111","0000110010001100100011001000","0000111111111111111111111111","0000111100101111001011110010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101111111011111110111","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000111110001111100011111000","0000111010101110101011101010","0000100010001000100010001000","0001000000000000000000000000","0000001001010010010100100101","0001000000000000000000000000","0000010001010100010101000101","0000100001101000011010000110","0000111010101110101011101010","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000110100011101000111010001","0000011010110110101101101011","0000100010011000100110001001","0000110100001101000011010000","0000011110110111101101111011","0001000000000000000000000000","0000000001010000010100000101","0000011010110110101101101011","0000111111111111111111111111","0000110111101101111011011110","0000110100111101001111010011","0000110110111101101111011011","0000111010001110100011101000","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111011111110111111101","0000111010011110100111101001","0000011101110111011101110111","0000110011101100111011001110","0000001111010011110100111101","0000110000011100000111000001",
		"0000111111111111111111111111","0000110011101100111011001110","0001000000000000000000000000","0000010111010101110101011101","0000101100101011001010110010","0000100111011001110110011101","0000110111001101110011011100","0000110100001101000011010000","0000111111001111110011111100","0000111110011111100111111001","0000111100101111001011110010","0000101000001010000010100000","0000110000011100000111000001","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111100011111000111110001","0000110011001100110011001100","0000111010101110101011101010","0000111011001110110011101100","0000100011001000110010001100","0000010010110100101101001011","0000001111010011110100111101","0000100100011001000110010001","0000101001111010011110100111","0000111110011111100111111001","0000011101000111010001110100","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110101111101011111010111","0000111000011110000111100001","0000011011000110110001101100","0000001111110011111100111111","0000110010111100101111001011","0000100011001000110010001100","0000111100011111000111110001","0000100111001001110010011100","0000100100011001000110010001","0000100010111000101110001011","0000111111111111111111111111","0000111100001111000011110000","0000111111001111110011111100","0000110101111101011111010111","0000110111111101111111011111","0000110111101101111011011110","0000111101111111011111110111","0000111111111111111111111111","0000111101001111010011110100","0000110111101101111011011110","0000100001101000011010000110","0000011011110110111101101111","0000010101000101010001010100","0000110100101101001011010010","0000011111110111111101111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111100111111001111110011","0000111101011111010111110101","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000101100011011000110110001","0000011101110111011101110111","0000011111010111110101111101","0000011011100110111001101110","0000011100110111001101110011","0000001100110011001100110011","0000011001100110011001100110","0000100100001001000010010000","0000010111100101111001011110","0000001111000011110000111100","0000001111110011111100111111","0000011000100110001001100010","0000000101000001010000010100","0001000000000000000000000000","0000100001001000010010000100","0000011101110111011101110111","0000010110000101100001011000","0000101100101011001010110010","0000111001001110010011100100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111111111111111111111111","0000111100101111001011110010","0000110110101101101011011010","0000100111001001110010011100","0000100101001001010010010100","0000011110010111100101111001","0000100011001000110010001100","0000011010110110101101101011","0000010001000100010001000100","0000000000110000001100000011","0000010001110100011101000111","0001000000000000000000000000","0000000011000000110000001100","0000000000010000000100000001","0000001100100011001000110010","0000101001101010011010100110","0000111100011111000111110001","0000111010011110100111101001","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110110001101100011011000","0000001100000011000000110000","0000010111100101111001011110","0000001110010011100100111001","0000001101110011011100110111","0000100010011000100110001001","0000111010001110100011101000","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111100111111001111110011","0000111100011111000111110001","0000111110001111100011111000","0000111000011110000111100001","0000101000111010001110100011","0000100010011000100110001001","0000101000101010001010100010","0000011001100110011001100110","0000001101000011010000110100","0000010100110101001101010011","0000101011011010110110101101","0000110100001101000011010000","0000100101101001011010010110","0000110111011101110111011101","0000111100101111001011110010","0000111101011111010111110101","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111110001111100011111000","0000111100011111000111110001","0000011100110111001101110011","0000101100101011001010110010","0000011000000110000001100000","0000100000101000001010000010",
		"0000111101001111010011110100","0000101001111010011110100111","0000000100000001000000010000","0000000101110001011100010111","0000100000111000001110000011","0000100000101000001010000010","0000101110111011101110111011","0000101111101011111010111110","0000111101011111010111110101","0000111111111111111111111111","0000101110101011101010111010","0000010010110100101101001011","0000111011001110110011101100","0000111111101111111011111110","0000111110001111100011111000","0000111100011111000111110001","0000111000101110001011100010","0000110011001100110011001100","0000111101011111010111110101","0000110001001100010011000100","0000100010001000100010001000","0000011101000111010001110100","0000001110100011101000111010","0000011111000111110001111100","0000101110101011101010111010","0000111000101110001011100010","0000101011101010111010101110","0000110011001100110011001100","0000111111101111111011111110","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111001101110011011100110","0000111111111111111111111111","0000110110001101100011011000","0000101011011010110110101101","0000100101011001010110010101","0000000011000000110000001100","0000011011010110110101101101","0000011110010111100101111001","0000100001101000011010000110","0000100010101000101010001010","0000011011110110111101101111","0000011100010111000101110001","0000101011111010111110101111","0000101011001010110010101100","0000101001001010010010100100","0000101100011011000110110001","0000110001011100010111000101","0000111001001110010011100100","0000111010111110101111101011","0000111111111111111111111111","0000111101011111010111110101","0000100100101001001010010010","0000100100101001001010010010","0000001111000011110000111100","0000011100000111000001110000","0000100101011001010110010101","0000110110111101101111011011","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111000111110001111100011","0000100110101001101010011010","0000101001101010011010100110","0000011011000110110001101100","0000011101010111010101110101","0000001000000010000000100000","0000010011000100110001001100","0000101001001010010010100100","0000010110100101101001011010","0000001110100011101000111010","0000001001100010011000100110","0000001011110010111100101111","0000000001010000010100000101","0000011011000110110001101100","0000011011000110110001101100","0000011100000111000001110000","0000110101011101010111010101","0000110011001100110011001100","0000100110111001101110011011","0000100110111001101110011011","0000101010111010101110101011","0000110000101100001011000010","0000110001001100010011000100","0000110101101101011011010110","0000110011001100110011001100","0000101110101011101010111010","0000101110111011101110111011","0000101010111010101110101011","0000100010101000101010001010","0000011010110110101101101011","0000010110010101100101011001","0000010011010100110101001101","0000010001010100010101000101","0000000111110001111100011111","0000000111000001110000011100","0000000110000001100000011000","0000000001000000010000000100","0000000011100000111000001110","0000000000100000001000000010","0000000010000000100000001000","0001000000000000000000000000","0000001010100010101000101010","0000010011100100111001001110","0000010000100100001001000010","0000011101100111011001110110","0000100001001000010010000100","0000101100001011000010110000","0000111001101110011011100110","0000110101101101011011010110","0000111001011110010111100101","0000111100101111001011110010","0000111111111111111111111111","0000111101101111011011110110","0000110110111101101111011011","0000111100011111000111110001","0000111111111111111111111111","0000111011001110110011101100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111110001111100011111000","0000111110001111100011111000","0000111111111111111111111111","0000111011111110111111101111","0000100011001000110010001100","0000001110000011100000111000","0000100001011000010110000101","0000001000010010000100100001","0000011111010111110101111101","0000111011011110110111101101","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000110111001101110011011100","0000101110111011101110111011","0000100010101000101010001010","0000011101100111011001110110","0000001001100010011000100110","0000000111010001110100011101","0000000001110000011100000111","0000011111110111111101111111","0000110001001100010011000100","0000110010011100100111001001","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111001111110011111100","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111001001110010011100100","0000100101011001010110010101","0000100111011001110110011101","0000011101000111010001110100","0000010010000100100001001000",
		"0000111110001111100011111000","0000011010000110100001101000","0000010101100101011001010110","0000010010110100101101001011","0000011101000111010001110100","0000011101000111010001110100","0000100100101001001010010010","0000100110111001101110011011","0000111111001111110011111100","0000110100011101000111010001","0000011001000110010001100100","0000110110111101101111011011","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000110110101101101011011010","0000110011111100111111001111","0000101011011010110110101101","0000010011100100111001001110","0000100100001001000010010000","0000000101000001010000010100","0000011111110111111101111111","0000100111011001110110011101","0000111111111111111111111111","0000111100111111001111110011","0000011101100111011001110110","0000111101011111010111110101","0000111110101111101011111010","0000111100001111000011110000","0000111110011111100111111001","0000111011101110111011101110","0000111111011111110111111101","0000111111111111111111111111","0000101110001011100010111000","0000100001111000011110000111","0000001001100010011000100110","0000000111110001111100011111","0000011001010110010101100101","0000010100100101001001010010","0000010100110101001101010011","0000010101110101011101010111","0000010000000100000001000000","0000011001000110010001100100","0000100010001000100010001000","0000101011101010111010101110","0000101110101011101010111010","0000110011001100110011001100","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000110110111101101111011011","0000100010101000101010001010","0000011111100111111001111110","0000010110000101100001011000","0000101010111010101110101011","0000100000011000000110000001","0000111101001111010011110100","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111010111110101111101011","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111010101110101011101010","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111011111110111111101","0000110101001101010011010100","0000111111001111110011111100","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111101001111010011110100","0000111110001111100011111000","0000111110101111101011111010","0000110110011101100111011001","0000100110011001100110011001","0000110001111100011111000111","0000010100110101001101010011","0000001010010010100100101001","0000000010110000101100001011","0000100110001001100010011000","0000100100101001001010010010","0000000010110000101100001011","0000000001000000010000000100","0000000010000000100000001000","0000000111000001110000011100","0000100001101000011010000110","0000010110100101101001011010","0000100101011001010110010101","0000111010101110101011101010","0000110001111100011111000111","0000101110101011101010111010","0000110000011100000111000001","0000100110101001101010011010","0000011011100110111001101110","0000010001010100010101000101","0000001111100011111000111110","0000001000010010000100100001","0000010001100100011001000110","0000010101000101010001010100","0000010110110101101101011011","0000010101100101011001010110","0000010111000101110001011100","0000011111000111110001111100","0000101001111010011110100111","0000110000111100001111000011","0000110111101101111011011110","0000110000111100001111000011","0000101000101010001010100010","0000100010111000101110001011","0000011001010110010101100101","0000011111100111111001111110","0000100101111001011110010111","0000101010111010101110101011","0000011101000111010001110100","0000011010110110101101101011","0000010110000101100001011000","0000100011011000110110001101","0000110001111100011111000111","0000101111101011111010111110","0000101110111011101110111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111100011111000111110001","0000111111111111111111111111","0000110010101100101011001010","0000101001011010010110100101","0000100100011001000110010001","0000100011111000111110001111","0000010111010101110101011101","0000111100111111001111110011","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111101001111010011110100","0000111111111111111111111111","0000110110001101100011011000","0000100001101000011010000110","0000011011010110110101101101","0000011100110111001101110011","0001000000000000000000000000","0001000000000000000000000000","0000011010010110100101101001","0000101111011011110110111101","0000100111111001111110011111","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111110101111101011111010","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111001111110011111100","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000110010011100100111001001","0000110001111100011111000111","0000100101011001010110010101","0000011100110111001101110011","0000001011110010111100101111",
		"0000111111111111111111111111","0000000101000001010000010100","0000010110110101101101011011","0000010110100101101001011010","0000001011000010110000101100","0000011011100110111001101110","0000100101101001011010010110","0000100011111000111110001111","0000100000101000001010000010","0000000100010001000100010001","0000110100111101001111010011","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111110001111100011111000","0000111010001110100011101000","0000110000101100001011000010","0000101011111010111110101111","0000100110111001101110011011","0000001100000011000000110000","0000011110000111100001111000","0001000000000000000000000000","0000100100111001001110010011","0000100000101000001010000010","0000111110001111100011111000","0000111111111111111111111111","0000101011101010111010101110","0000100111011001110110011101","0000110100111101001111010011","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000110010101100101011001010","0000100000001000000010000000","0001000000000000000000000000","0000010000000100000001000000","0000011000110110001101100011","0000010001010100010101000101","0000010111100101111001011110","0000011100010111000101110001","0000011101000111010001110100","0000110000111100001111000011","0000111111111111111111111111","0000111010011110100111101001","0000111110011111100111111001","0000111011001110110011101100","0000111101111111011111110111","0000111111111111111111111111","0000101100001011000010110000","0000100000001000000010000000","0000011111100111111001111110","0000100010001000100010001000","0000101010111010101110101011","0000101110111011101110111011","0000110111111101111111011111","0000110100101101001011010010","0000111110111111101111111011","0000111111101111111011111110","0000111100111111001111110011","0000111101001111010011110100","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111010101110101011101010","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000110110011101100111011001","0000110010111100101111001011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000110100001101000011010000","0000110110001101100011011000","0000100001001000010010000100","0000100000011000000110000001","0000000110010001100100011001","0000010001000100010001000100","0000100001001000010010000100","0001000000000000000000000000","0000000001110000011100000111","0000001010100010101000101010","0000001001110010011100100111","0000100110001001100010011000","0000010110010101100101011001","0000011001010110010101100101","0000111101011111010111110101","0000111100101111001011110010","0000101010101010101010101010","0000010100110101001101010011","0000001111000011110000111100","0000001111010011110100111101","0000011010010110100101101001","0000011101010111010101110101","0000011101000111010001110100","0000100101101001011010010110","0000101110001011100010111000","0000110110011101100111011001","0000111000101110001011100010","0000110111111101111111011111","0000110111111101111111011111","0000111000111110001111100011","0000111000111110001111100011","0000110101111101011111010111","0000110011011100110111001101","0000110001111100011111000111","0000101111101011111010111110","0000011100000111000001110000","0000011111100111111001111110","0000011100100111001001110010","0000011100000111000001110000","0000100010001000100010001000","0000100111111001111110011111","0000011110100111101001111010","0000100010011000100110001001","0000110001111100011111000111","0000111100111111001111110011","0000111111111111111111111111","0000111011101110111011101110","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111101101111011011110110","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111100101111001011110010","0000111110111111101111111011","0000110011011100110111001101","0000100010011000100110001001","0000100110111001101110011011","0000011101000111010001110100","0000111001001110010011100100","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111101001111010011110100","0000111111111111111111111111","0000111111001111110011111100","0000110110101101101011011010","0000101011001010110010101100","0000100100011001000110010001","0000011110100111101001111010","0000010001000100010001000100","0000000011000000110000001100","0000001010010010100100101001","0000101110111011101110111011","0000101001101010011010100110","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111011111110111111101","0000111110111111101111111011","0000101100001011000010110000","0000110110111101101111011011","0000100101011001010110010101","0000010110000101100001011000","0000001110010011100100111001",
		"0000111000011110000111100001","0000000100100001001000010010","0000101001101010011010100110","0000100000111000001110000011","0000000101110001011100010111","0000001110010011100100111001","0000001110100011101000111010","0001000000000000000000000000","0000000000100000001000000010","0000101110011011100110111001","0000111111001111110011111100","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111000001110000011100000","0000101000111010001110100011","0000100110101001101010011010","0000100001101000011010000110","0000000101100001011000010110","0000100001101000011010000110","0000000110100001101000011010","0000100100101001001010010010","0000011111100111111001111110","0000110100101101001011010010","0000111010011110100111101001","0000111111111111111111111111","0000110000011100000111000001","0000010110010101100101011001","0000111011111110111111101111","0000111010101110101011101010","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000110010111100101111001011","0000010010100100101001001010","0000001001100010011000100110","0000010010100100101001001010","0000010101010101010101010101","0000010000100100001001000010","0000100110111001101110011011","0000011010000110100001101000","0000101110001011100010111000","0000111000101110001011100010","0000111010101110101011101010","0000111011111110111111101111","0000111101011111010111110101","0000110010001100100011001000","0000111110011111100111111001","0000101000101010001010100010","0000010111110101111101011111","0000101000001010000010100000","0000011110000111100001111000","0000101001011010010110100101","0000101000111010001110100011","0000111111111111111111111111","0000100111011001110110011101","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111101001111010011110100","0000111011011110110111101101","0000111011111110111111101111","0000111011111110111111101111","0000111011001110110011101100","0000111100101111001011110010","0000111111101111111011111110","0000111110111111101111111011","0000111000101110001011100010","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111100001111000011110000","0000101100001011000010110000","0000111100001111000011110000","0000111100101111001011110010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111101001111010011110100","0000101110011011100110111001","0000101001101010011010100110","0000011001100110011001100110","0000010001010100010101000101","0000000101110001011100010111","0000001111010011110100111101","0000001010110010101100101011","0000000010010000100100001001","0000001000010010000100100001","0000000010010000100100001001","0000100100001001000010010000","0000101110101011101010111010","0000001110110011101100111011","0000101000001010000010100000","0000100001111000011110000111","0000011000110110001101100011","0000011010000110100001101000","0000110001001100010011000100","0000111001111110011111100111","0000110100111101001111010011","0000110000101100001011000010","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111011001110110011101100","0000111100101111001011110010","0000111101101111011011110110","0000111101011111010111110101","0000111111111111111111111111","0000111110001111100011111000","0000111011101110111011101110","0000110011101100111011001110","0000100011111000111110001111","0000101001011010010110100101","0000101000011010000110100001","0000101001001010010010100100","0000110000001100000011000000","0000101111111011111110111111","0000111111111111111111111111","0000111011011110110111101101","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110111101101111011011110","0000110110011101100111011001","0000111111101111111011111110","0000111101111111011111110111","0000111010001110100011101000","0000111111011111110111111101","0000111111001111110011111100","0000111011011110110111101101","0000111110011111100111111001","0000111101111111011111110111","0000111011111110111111101111","0000111101011111010111110101","0000111001111110011111100111","0000100010111000101110001011","0000011001110110011101100111","0000011010000110100001101000","0000101000101010001010100010","0000111111001111110011111100","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000110101001101010011010100","0000101011101010111010101110","0000011110110111101101111011","0000010000000100000001000000","0000001100100011001000110010","0000001100110011001100110011","0000011110010111100101111001","0000101110111011101110111011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011111110111111101111","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111011111110111111101","0000101001101010011010100110","0000110000111100001111000011","0000100110001001100010011000","0000001010010010100100101001","0000010010110100101101001011",
		"0000110011011100110111001101","0001000000000000000000000000","0000101101101011011010110110","0000101110001011100010111000","0000010110100101101001011010","0000000010010000100100001001","0000001110100011101000111010","0000100010101000101010001010","0000110000111100001111000011","0000111011011110110111101101","0000111100011111000111110001","0000111110001111100011111000","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111100001111000011110000","0000111100101111001011110010","0000011001000110010001100100","0000011100100111001001110010","0000100010111000101110001011","0000001100110011001100110011","0000100000111000001110000011","0000001100000011000000110000","0000101001011010010110100101","0000011100000111000001110000","0000101111101011111010111110","0000111111111111111111111111","0000111001101110011011100110","0000110111101101111011011110","0000100010111000101110001011","0000101101011011010110110101","0000101001001010010010100100","0000101001011010010110100101","0000101110011011100110111001","0000101010111010101110101011","0000100111111001111110011111","0000100101111001011110010111","0000010111100101111001011110","0000011100010111000101110001","0001000000000000000000000000","0000001100000011000000110000","0000010011000100110001001100","0000010100110101001101010011","0000010000110100001101000011","0000011101010111010101110101","0000001010100010101000101010","0000101001011010010110100101","0000110011011100110111001101","0000110001001100010011000100","0000110111001101110011011100","0000111111011111110111111101","0000100111001001110010011100","0000100101011001010110010101","0000101000101010001010100010","0000011001110110011101100111","0000011001000110010001100100","0000101001001010010010100100","0000100101011001010110010101","0000111000011110000111100001","0000110000011100000111000001","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000110101111101011111010111","0000110100101101001011010010","0000111010101110101011101010","0000111111111111111111111111","0000111110011111100111111001","0000111000011110000111100001","0000111000001110000011100000","0000111111111111111111111111","0000111001011110010111100101","0000111101101111011011110110","0000111111111111111111111111","0000111001001110010011100100","0000110101011101010111010101","0000101111001011110010111100","0000111111011111110111111101","0000111110111111101111111011","0000111110011111100111111001","0000111101111111011111110111","0000111101011111010111110101","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000101111111011111110111111","0000000110010001100100011001","0000100111001001110010011100","0000010010100100101001001010","0000000000110000001100000011","0000000101000001010000010100","0000000100000001000000010000","0001000000000000000000000000","0000000001000000010000000100","0000010110100101101001011010","0000110111011101110111011101","0000010011000100110001001100","0000011000010110000101100001","0000011001110110011101100111","0000100011111000111110001111","0000101100001011000010110000","0000101101101011011010110110","0000110111011101110111011101","0000111000101110001011100010","0000111100101111001011110010","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111101101111011011110110","0000111111111111111111111111","0000111111001111110011111100","0000111010001110100011101000","0000111100111111001111110011","0000111101101111011011110110","0000111100011111000111110001","0000110010111100101111001011","0000101100001011000010110000","0000110000011100000111000001","0000110010101100101011001010","0000101101101011011010110110","0000101001111010011110100111","0000100001001000010010000100","0000111011011110110111101101","0000111011111110111111101111","0000110011101100111011001110","0000111111101111111011111110","0000111111111111111111111111","0000111010011110100111101001","0000111110011111100111111001","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000111100111111001111110011","0000110101101101011011010110","0000010110000101100001011000","0000101000011010000110100001","0000101111101011111010111110","0000111111001111110011111100","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111101011111010111110101","0000111111001111110011111100","0000111100001111000011110000","0000101001011010010110100101","0000100011001000110010001100","0000011100110111001101110011","0000001110110011101100111011","0000011000100110001001100010","0000011001100110011001100110","0000110010111100101111001011","0000111111011111110111111101","0000111110011111100111111001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111110111111101111111011","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110001111100011111000","0000111101101111011011110110","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111101111111011111110111","0000111111011111110111111101","0000101001011010010110100101","0000101000011010000110100001","0000100110101001101010011010","0000000000010000000100000001","0000010101000101010001010100",
		"0000101101111011011110110111","0000010100110101001101010011","0000101000001010000010100000","0000110110101101101011011010","0000011111110111111101111111","0001000000000000000000000000","0000011011110110111101101111","0000011111010111110101111101","0000111010111110101111101011","0000111101101111011011110110","0000111100101111001011110010","0000111111001111110011111100","0000111101111111011111110111","0000111101001111010011110100","0000111111111111111111111111","0000111101011111010111110101","0000111100101111001011110010","0000010110110101101101011011","0000010010010100100101001001","0000011101100111011001110110","0000010101110101011101010111","0000011000110110001101100011","0000011010110110101101101011","0000011010010110100101101001","0000100010011000100110001001","0000110001111100011111000111","0000111111111111111111111111","0000110110001101100011011000","0000111001101110011011100110","0000011110100111101001111010","0000101110101011101010111010","0000101000101010001010100010","0000101011001010110010101100","0000011001100110011001100110","0000000110010001100100011001","0000001001100010011000100110","0000010010000100100001001000","0000010011100100111001001110","0000010110110101101101011011","0000010101000101010001010100","0000001111100011111000111110","0000000100110001001100010011","0001000000000000000000000000","0000001110000011100000111000","0000010100010101000101010001","0000010111000101110001011100","0000100001111000011110000111","0000101110011011100110111001","0000111111111111111111111111","0000111100001111000011110000","0000110000111100001111000011","0000100111111001111110011111","0000100011111000111110001111","0000101011111010111110101111","0000011111110111111101111111","0000011101010111010101110101","0000010110000101100001011000","0000100010101000101010001010","0000111110011111100111111001","0000101010011010100110101001","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000110110101101101011011010","0000110011101100111011001110","0000110100101101001011010010","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000101111001011110010111100","0000111110001111100011111000","0000111111011111110111111101","0000111100111111001111110011","0000111110011111100111111001","0000111111011111110111111101","0000111011011110110111101101","0000111101101111011011110110","0000111110011111100111111001","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000110000101100001011000010","0000101000011010000110100001","0000110110011101100111011001","0000011110110111101101111011","0000000011010000110100001101","0000000010010000100100001001","0000001100110011001100110011","0001000000000000000000000000","0000010101100101011001010110","0000011111000111110001111100","0000100011001000110010001100","0000010100010101000101010001","0000100001111000011110000111","0000101001101010011010100110","0000010100100101001001010010","0000011111010111110101111101","0000100101111001011110010111","0000101111111011111110111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111100101111001011110010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000111000011110000111100001","0000111101011111010111110101","0000111111111111111111111111","0000111010101110101011101010","0000111011011110110111101101","0000110000011100000111000001","0000110011011100110111001101","0000100011101000111010001110","0000011011000110110001101100","0000100011011000110110001101","0000110110101101101011011010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111101111111011111110111","0000111101001111010011110100","0000111101001111010011110100","0000111110111111101111111011","0000111010001110100011101000","0000101101001011010010110100","0000101010101010101010101010","0000111000001110000011100000","0000110101011101010111010101","0000111101111111011111110111","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000110110011101100111011001","0000101101001011010010110100","0000110100111101001111010011","0000101111001011110010111100","0000110000001100000011000000","0000011011110110111101101111","0000000101000001010000010100","0000010011110100111101001111","0000110010101100101011001010","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111110101111101011111010","0000111111101111111011111110","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000110110101101101011011010","0000111111111111111111111111","0000111101011111010111110101","0000111111001111110011111100","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000110001011100010111000101","0000101100101011001010110010","0000101001101010011010100110","0001000000000000000000000000","0000011100110111001101110011",
		"0000100101101001011010010110","0000010000100100001001000010","0000110100111101001111010011","0000110010101100101011001010","0000010111110101111101011111","0000011100010111000101110001","0000001000010010000100100001","0000101101101011011010110110","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111100111111001111110011","0000111111111111111111111111","0000111100101111001011110010","0000111110111111101111111011","0000111111111111111111111111","0000101010001010100010101000","0000011000000110000001100000","0000010011110100111101001111","0000100000001000000010000000","0000000111110001111100011111","0000100111111001111110011111","0000101011001010110010101100","0000001111000011110000111100","0000100011111000111110001111","0000110000001100000011000000","0000111100001111000011110000","0000110011101100111011001110","0000110101111101011111010111","0000100101101001011010010110","0000110000101100001011000010","0000100010101000101010001010","0000010001010100010101000101","0000010010100100101001001010","0000010011110100111101001111","0000011000110110001101100011","0000011101010111010101110101","0000100010001000100010001000","0000101011011010110110101101","0000110001001100010011000100","0000110001011100010111000101","0000111000001110000011100000","0000101111011011110110111101","0000011100100111001001110010","0000000001000000010000000100","0000001100100011001000110010","0000010101110101011101010111","0000001000110010001100100011","0000001101110011011100110111","0000010011110100111101001111","0000100000001000000010000000","0000100111011001110110011101","0000100100101001001010010010","0000011000000110000001100000","0000011111100111111001111110","0000011101100111011001110110","0000010100010101000101010001","0000010110000101100001011000","0000110111111101111111011111","0000100110101001101010011010","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111001101110011011100110","0000111000101110001011100010","0000111011001110110011101100","0000110011101100111011001110","0000101101101011011010110110","0000101011011010110110101101","0000110000011100000111000001","0000101110111011101110111011","0000110010111100101111001011","0000110111111101111111011111","0000111101001111010011110100","0000111100101111001011110010","0000111101001111010011110100","0000101100111011001110110011","0000111111111111111111111111","0000111101101111011011110110","0000111011101110111011101110","0000111101101111011011110110","0000111001101110011011100110","0000111101011111010111110101","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111010101110101011101010","0000100100111001001110010011","0000111010001110100011101000","0000100001101000011010000110","0001000000000000000000000000","0000000010100000101000001010","0000001010110010101100101011","0000000100000001000000010000","0000001101010011010100110101","0000011110100111101001111010","0000100010101000101010001010","0000010100010101000101010001","0000110010101100101011001010","0000101100111011001110110011","0000100010111000101110001011","0000101100001011000010110000","0000110111111101111111011111","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111111101111111011111110","0000111100011111000111110001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111101101111011011110110","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000110101111101011111010111","0000101100111011001110110011","0000100001101000011010000110","0000100101001001010010010100","0000010110000101100001011000","0000010111010101110101011101","0000110000001100000011000000","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000110010001100100011001000","0000110001011100010111000101","0000100110011001100110011001","0000111100001111000011110000","0000111111011111110111111101","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111001101110011011100110","0000101011111010111110101111","0000101001001010010010100100","0000110011011100110111001101","0000101100011011000110110001","0000111110101111101011111010","0000011110000111100001111000","0000011001110110011101100111","0000000011110000111100001111","0000100100101001001010010010","0000111000101110001011100010","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000110111111101111111011111","0000111000011110000111100001","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111101011111010111110101","0000101100111011001110110011","0000101110101011101010111010","0000101100001011000010110000","0000001000100010001000100010","0000100100001001000010010000",
		"0000011001110110011101100111","0000011000110110001101100011","0000110101011101010111010101","0000101001011010010110100101","0000011100010111000101110001","0000011110010111100101111001","0000001011000010110000101100","0000110101001101010011010100","0000111011011110110111101101","0000111101111111011111110111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000110000101100001011000010","0000011011000110110001101100","0000011000010110000101100001","0000010101100101011001010110","0000010101100101011001010110","0000010010100100101001001010","0000110100011101000111010001","0000111001111110011111100111","0000000011100000111000001110","0000100101111001011110010111","0000101110001011100010111000","0000111100011111000111110001","0000110110001101100011011000","0000111010011110100111101001","0000101000001010000010100000","0000111111111111111111111111","0000111010111110101111101011","0000111011011110110111101101","0000111100111111001111110011","0000111110011111100111111001","0000111010011110100111101001","0000111000101110001011100010","0000111011011110110111101101","0000111100101111001011110010","0000111110101111101011111010","0000111111001111110011111100","0000110111101101111011011110","0000111010111110101111101011","0000111001001110010011100100","0000110011001100110011001100","0000011001100110011001100110","0000011001110110011101100111","0000011011110110111101101111","0000100100011001000110010001","0000101010101010101010101010","0000100001011000010110000101","0000011001010110010101100101","0000010001010100010101000101","0000001101110011011100110111","0000010011010100110101001101","0000010100100101001001010010","0000011000110110001101100011","0000010000000100000001000000","0000101010001010100010101000","0000101011001010110010101100","0000101100101011001010110010","0000111011101110111011101110","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000110111111101111111011111","0000101011001010110010101100","0000100000011000000110000001","0000100000001000000010000000","0000100011001000110010001100","0000101001111010011110100111","0000110000101100001011000010","0000110100101101001011010010","0000110110001101100011011000","0000110010011100100111001001","0000111011001110110011101100","0000110110001101100011011000","0000110111111101111111011111","0000111001001110010011100100","0000111111111111111111111111","0000101100101011001010110010","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111010001110100011101000","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000101111111011111110111111","0000111100101111001011110010","0000101111101011111010111110","0000000011110000111100001111","0000000101000001010000010100","0000001111000011110000111100","0000000011010000110100001101","0000000000110000001100000011","0000100011101000111010001110","0000010111000101110001011100","0000011100010111000101110001","0000110110001101100011011000","0000100010001000100010001000","0000101100111011001110110011","0000101100101011001010110010","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111110011111100111111001","0000111110101111101011111010","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111010111110101111101011","0000111010111110101111101011","0000111001111110011111100111","0000101100011011000110110001","0000010011000100110001001100","0000010001100100011001000110","0000100001101000011010000110","0000111010011110100111101001","0000111101111111011111110111","0000111110001111100011111000","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000101011011010110110101101","0000111011101110111011101110","0000110001101100011011000110","0000110001101100011011000110","0000111101001111010011110100","0000111111111111111111111111","0000111110001111100011111000","0000111000101110001011100010","0000101101101011011010110110","0000110100111101001111010011","0000110101011101010111010101","0000111100101111001011110010","0000101111111011111110111111","0000111111111111111111111111","0000001111000011110000111100","0000100101101001011010010110","0000000100000001000000010000","0000011000000110000001100000","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111100001111000011110000","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000110011011100110111001101","0000111001101110011011100110","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111110111111101111111011","0000111111111111111111111111","0000101111111011111110111111","0000101111111011111110111111","0000100001101000011010000110","0001000000000000000000000000","0000101100011011000110110001",
		"0000010100000101000001010000","0000101011101010111010101110","0000110010001100100011001000","0000101010001010100010101000","0000100010111000101110001011","0000010010100100101001001010","0000100010101000101010001010","0000111011001110110011101100","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111110101111101011111010","0000101111101011111010111110","0000100001101000011010000110","0000100101011001010110010101","0000101010011010100110101001","0000000110100001101000011010","0000000111010001110100011101","0000011111110111111101111111","0000111100011111000111110001","0000110100101101001011010010","0000010010110100101101001011","0000100000101000001010000010","0000101100011011000110110001","0000110001111100011111000111","0000110010101100101011001010","0000111001101110011011100110","0000101100011011000110110001","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000110100011101000111010001","0000101101111011011110110111","0000110001001100010011000100","0000101100111011001110110011","0000101011101010111010101110","0000100111001001110010011100","0000011111000111110001111100","0000011010010110100101101001","0000100000111000001110000011","0000101011001010110010101100","0000101111011011110110111101","0000110111111101111111011111","0000100001001000010010000100","0000011000110110001101100011","0000001001110010011100100111","0000001001100010011000100110","0000001110110011101100111011","0000100010101000101010001010","0000011010010110100101101001","0000010010110100101101001011","0000101011001010110010101100","0000100101011001010110010101","0000100111101001111010011110","0000101011011010110110101101","0000110000001100000011000000","0000101111101011111010111110","0000101111001011110010111100","0000101011101010111010101110","0000100011001000110010001100","0000011100110111001101110011","0000011010100110101001101010","0000011001000110010001100100","0000011000010110000101100001","0000011111000111110001111100","0000011100110111001101110011","0000011101010111010101110101","0000011010110110101101101011","0000100011001000110010001100","0000100110101001101010011010","0000110100101101001011010010","0000110011001100110011001100","0000101111111011111110111111","0000110101011101010111010101","0000111111111111111111111111","0000111111001111110011111100","0000111011101110111011101110","0000111111001111110011111100","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111011101110111011101110","0000100011101000111010001110","0000111001101110011011100110","0000101111011011110110111101","0000010111100101111001011110","0001000000000000000000000000","0000010010010100100101001001","0000000111010001110100011101","0000000010010000100100001001","0000011001010110010101100101","0000001011010010110100101101","0000011010110110101101101011","0000110110011101100111011001","0000101010001010100010101000","0000110010111100101111001011","0000110010111100101111001011","0000111101111111011111110111","0000111010101110101011101010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110111111101111111011","0000111011101110111011101110","0000111011111110111111101111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111101101111011011110110","0000110111011101110111011101","0000111111111111111111111111","0000110010111100101111001011","0000010110100101101001011010","0000010011010100110101001101","0000011100010111000101110001","0000101101001011010010110100","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111100101111001011110010","0000111110101111101011111010","0000111110101111101011111010","0000111100111111001111110011","0000101000001010000010100000","0000111111111111111111111111","0000111111111111111111111111","0000110101111101011111010111","0000111101101111011011110110","0000111100101111001011110010","0000111011001110110011101100","0000101000101010001010100010","0000100111001001110010011100","0000111111101111111011111110","0000110111011101110111011101","0000111000111110001111100011","0000110111011101110111011101","0000011111100111111001111110","0000100111101001111010011110","0000011110110111101101111011","0000001010010010100100101001","0000101001101010011010100110","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111100011111000111110001","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000110101011101010111010101","0000111001011110010111100101","0000110110001101100011011000","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111101011111010111110101","0000101001011010010110100101","0000110001011100010111000101","0000100010011000100110001001","0001000000000000000000000000","0000110100111101001111010011",
		"0000000111100001111000011110","0000101110111011101110111011","0000110110001101100011011000","0000101110001011100010111000","0000010011000100110001001100","0000010001010100010101000101","0000101000101010001010100010","0000111111001111110011111100","0000111100011111000111110001","0000111111111111111111111111","0000111001111110011111100111","0000111100111111001111110011","0000111101101111011011110110","0000110100101101001011010010","0000100001111000011110000111","0000100100011001000110010001","0000101001101010011010100110","0000001101010011010100110101","0000000010110000101100001011","0000100010011000100110001001","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000011000100110001001100010","0000001001000010010000100100","0000100111011001110110011101","0000101101001011010010110100","0000110001001100010011000100","0000110011001100110011001100","0000110010111100101111001011","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111110011111100111111001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110111001101110011011100","0000111000101110001011100010","0000101100001011000010110000","0000101110001011100010111000","0000100110101001101010011010","0000110000011100000111000001","0000101100101011001010110010","0000101101101011011010110110","0000100001001000010010000100","0000100011011000110110001101","0000101011001010110010101100","0000010011000100110001001100","0000001110100011101000111010","0000000101110001011100010111","0000001011100010111000101110","0000010100010101000101010001","0000100011001000110010001100","0000001011100010111000101110","0000010101000101010001010100","0000011100110111001101110011","0000100000011000000110000001","0000011110100111101001111010","0000011001000110010001100100","0000011110110111101101111011","0000010110100101101001011010","0000001000010010000100100001","0001000000000000000000000000","0001000000000000000000000000","0000000001110000011100000111","0000000110110001101100011011","0000000111000001110000011100","0001000000000000000000000000","0000000010010000100100001001","0000000101000001010000010100","0000001110100011101000111010","0000010001000100010001000100","0000011110010111100101111001","0000100101011001010110010101","0000110110111101101111011011","0000101110111011101110111011","0000101111111011111110111111","0000111001101110011011100110","0000110111101101111011011110","0000101010011010100110101001","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110001111100011111000","0000111110111111101111111011","0000111110001111100011111000","0000111111011111110111111101","0000101101101011011010110110","0000111100101111001011110010","0000101110011011100110111001","0000101010001010100010101000","0000000011000000110000001100","0000001000100010001000100010","0000000111100001111000011110","0000000110000001100000011000","0000010000000100000001000000","0000010111000101110001011100","0000010101010101010101010101","0000110010111100101111001011","0000110011111100111111001111","0000100110111001101110011011","0000111010011110100111101001","0000111011101110111011101110","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111010011110100111101001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000110011111100111111001111","0000111110011111100111111001","0000101110101011101010111010","0000010101110101011101010111","0000011000100110001001100010","0000100101011001010110010101","0000100000111000001110000011","0000111011111110111111101111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111011101110111011101110","0000110101101101011011010110","0000111111111111111111111111","0000111100111111001111110011","0000111100011111000111110001","0000111110001111100011111000","0000110111001101110011011100","0000101000001010000010100000","0000100001101000011010000110","0000111110111111101111111011","0000110001101100011011000110","0000111110111111101111111011","0000111001011110010111100101","0000011110110111101101111011","0000100001001000010010000100","0000011001110110011101100111","0000001111010011110100111101","0000100011001000110010001100","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111011001110110011101100","0000111111101111111011111110","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000110010111100101111001011","0000111011101110111011101110","0000101011101010111010101110","0000111011111110111111101111","0000111111101111111011111110","0000111101101111011011110110","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110011001100110011001100","0000101111101011111010111110","0000001111010011110100111101","0000010111100101111001011110","0000111111111111111111111111",
		"0001000000000000000000000000","0000101101101011011010110110","0000111111111111111111111111","0000101101111011011110110111","0000001011000010110000101100","0000010000110100001101000011","0000101000011010000110100001","0000111110111111101111111011","0000111110111111101111111011","0000110010111100101111001011","0000111100011111000111110001","0000111111011111110111111101","0000110100001101000011010000","0000101111011011110110111101","0000101011101010111010101110","0000011111000111110001111100","0000000000110000001100000011","0000001010010010100100101001","0000100101001001010010010100","0000101100001011000010110000","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000011010010110100101101001","0000000100010001000100010001","0000011000010110000101100001","0000110010011100100111001001","0000101001101010011010100110","0000110010111100101111001011","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000110110001101100011011000","0000101111011011110110111101","0000101101001011010010110100","0000110001011100010111000101","0000110101101101011011010110","0000110100111101001111010011","0000110001011100010111000101","0000110001001100010011000100","0000101111101011111010111110","0000110000111100001111000011","0000100100101001001010010010","0000011111000111110001111100","0000010111110101111101011111","0000100001001000010010000100","0000010001000100010001000100","0000000111010001110100011101","0000001111010011110100111101","0000001101110011011100110111","0000010001100100011001000110","0000011001010110010101100101","0000011000010110000101100001","0000011110010111100101111001","0000100000001000000010000000","0000010110100101101001011010","0000010001000100010001000100","0000010010100100101001001010","0000010111000101110001011100","0000001100010011000100110001","0000001000010010000100100001","0001000000000000000000000000","0001000000000000000000000000","0000001101110011011100110111","0000100010011000100110001001","0000101010001010100010101000","0000101010001010100010101000","0000100101101001011010010110","0000100010101000101010001010","0000010110100101101001011010","0000001100010011000100110001","0000000110110001101100011011","0000000000110000001100000011","0000000111100001111000011110","0000010010110100101101001011","0000101111001011110010111100","0000100000011000000110000001","0000100001001000010010000100","0000111010101110101011101010","0000110011101100111011001110","0000101011001010110010101100","0000111011111110111111101111","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000110111111101111111011111","0000110110111101101111011011","0000111010001110100011101000","0000110011101100111011001110","0000111010111110101111101011","0000010000110100001101000011","0001000000000000000000000000","0000000101000001010000010100","0000000001000000010000000100","0000011101010111010101110101","0000011000110110001101100011","0000011101000111010001110100","0000101001111010011110100111","0000101101011011010110110101","0000011110110111101101111011","0000111001011110010111100101","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111000011110000111100001","0000111010011110100111101001","0000111011101110111011101110","0000110111001101110011011100","0000111111111111111111111111","0000111110011111100111111001","0000101111001011110010111100","0000110100101101001011010010","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000101101101011011010110110","0000111110111111101111111011","0000111110111111101111111011","0000100100111001001110010011","0000001101110011011100110111","0000100110001001100010011000","0000101011101010111010101110","0000100011111000111110001111","0000110100001101000011010000","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011011110110111101101","0000111111101111111011111110","0000111101011111010111110101","0000111011001110110011101100","0000111100001111000011110000","0000111101001111010011110100","0000101001001010010010100100","0000011101010111010101110101","0000111001011110010111100101","0000101011111010111110101111","0000111011111110111111101111","0000111010111110101111101011","0000110000011100000111000001","0000101011001010110010101100","0000011001100110011001100110","0001000000000000000000000000","0000110010011100100111001001","0000110001101100011011000110","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000110111011101110111011101","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000110011001100110011001100","0000110011111100111111001111","0000011110100111101001111010","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000001110000011100000","0000110000111100001111000011","0000101110101011101010111010","0000001110100011101000111010","0000011011010110110101101101","0000111111111111111111111111",
		"0000001000000010000000100000","0000110101111101011111010111","0000111111111111111111111111","0000101010011010100110101001","0000010111100101111001011110","0000001101010011010100110101","0000100111101001111010011110","0000111110001111100011111000","0000101011101010111010101110","0000111000111110001111100011","0000101111101011111010111110","0000101110011011100110111001","0000101010011010100110101001","0000110000111100001111000011","0000011101000111010001110100","0000100010011000100110001001","0000101111101011111010111110","0000100000001000000010000000","0000101100011011000110110001","0000111101001111010011110100","0000111110111111101111111011","0000111110011111100111111001","0000111110011111100111111001","0000101110111011101110111011","0000010111000101110001011100","0000000101100001011000010110","0000101110101011101010111010","0000011100100111001001110010","0000101100011011000110110001","0000100110011001100110011001","0000110100111101001111010011","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111101011111010111110101","0000111101011111010111110101","0000111110011111100111111001","0000111011111110111111101111","0000110100001101000011010000","0000110101101101011011010110","0000110100001101000011010000","0000110000101100001011000010","0000110101001101010011010100","0000100111011001110110011101","0000011001100110011001100110","0000100010001000100010001000","0000010111010101110101011101","0000010111110101111101011111","0000010010010100100101001001","0000010110000101100001011000","0000010111000101110001011100","0000101100011011000110110001","0000101100001011000010110000","0000001101010011010100110101","0000010000100100001001000010","0001000000000000000000000000","0000010011010100110101001101","0000010101010101010101010101","0000000011110000111100001111","0000000001100000011000000110","0000010001000100010001000100","0000011011000110110001101100","0000100011111000111110001111","0000110100011101000111010001","0000111100111111001111110011","0000111100011111000111110001","0000110011111100111111001111","0000101011101010111010101110","0000101000111010001110100011","0000100010101000101010001010","0000011111110111111101111111","0000010110000101100001011000","0000010101010101010101010101","0000010101000101010001010100","0000010011100100111001001110","0000001100110011001100110011","0000001000110010001100100011","0000000101010001010100010101","0000011011000110110001101100","0000011100100111001001110010","0000011011100110111001101110","0000101101001011010010110100","0000100110101001101010011010","0000110110111101101111011011","0000111101111111011111110111","0000111111111111111111111111","0000111011011110110111101101","0000111111001111110011111100","0000111100011111000111110001","0000111101011111010111110101","0000110111111101111111011111","0000111010001110100011101000","0000101010101010101010101010","0000101110101011101010111010","0000100000101000001010000010","0001000000000000000000000000","0000001111000011110000111100","0001000000000000000000000000","0000101000011010000110100001","0000000100110001001100010011","0000011011000110110001101100","0000100110011001100110011001","0000101111011011110110111101","0000101100101011001010110010","0000110111111101111111011111","0000111111111111111111111111","0000111100001111000011110000","0000111010011110100111101001","0000101110101011101010111010","0000110000101100001011000010","0000111000011110000111100001","0000111101101111011011110110","0000101101011011010110110101","0000101001001010010010100100","0000111111101111111011111110","0000111111111111111111111111","0000110111011101110111011101","0000111100001111000011110000","0000111011111110111111101111","0000111100001111000011110000","0000111100111111001111110011","0000111101011111010111110101","0000111110001111100011111000","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111100011111000111110001","0000100110101001101010011010","0000111100001111000011110000","0000101110111011101110111011","0000011110110111101101111011","0000010000110100001101000011","0000110100011101000111010001","0000101101111011011110110111","0000100110001001100010011000","0000110001001100010011000100","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111101101111011011110110","0000111011111110111111101111","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000101100011011000110110001","0000010110100101101001011010","0000101101011011010110110101","0000101100111011001110110011","0000110011011100110111001101","0000111101111111011111110111","0000101111011011110110111101","0000111111111111111111111111","0000011110000111100001111000","0001000000000000000000000000","0000101010001010100010101000","0000111001001110010011100100","0000110100101101001011010010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110101111101011111010111","0000111111011111110111111101","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000111000001110000011100000","0000101011111010111110101111","0000010110110101101101011011","0000110100011101000111010001","0000111100101111001011110010","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000110110111101101111011011","0000111001111110011111100111","0000101100101011001010110010","0000000010010000100100001001","0000010111100101111001011110","0000111000011110000111100001",
		"0000010100000101000001010000","0000110110111101101111011011","0000110101111101011111010111","0000100000111000001110000011","0000011010100110101001101010","0000001000100010001000100010","0000010111110101111101011111","0000111000001110000011100000","0000110000111100001111000011","0000101001001010010010100100","0000110110001101100011011000","0000101000101010001010100010","0000110011101100111011001110","0000110011011100110111001101","0000111111111111111111111111","0000111100111111001111110011","0000111010101110101011101010","0000101110111011101110111011","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111101011111010111110101","0000111111111111111111111111","0000110101101101011011010110","0000010111010101110101011101","0001000000000000000000000000","0000101111001011110010111100","0000100001001000010010000100","0000011110100111101001111010","0000101100101011001010110010","0000101101111011011110110111","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000101110111011101110111011","0000101001001010010010100100","0000100010001000100010001000","0000011100100111001001110010","0000100001111000011110000111","0000100101111001011110010111","0000110001101100011011000110","0000101011101010111010101110","0000101110111011101110111011","0000100111101001111010011110","0000100001111000011110000111","0000100100011001000110010001","0000100011111000111110001111","0000111001001110010011100100","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000101101101011011010110110","0000101101011011010110110101","0000101110101011101010111010","0000100010111000101110001011","0000011000110110001101100011","0000101000111010001110100011","0000101111011011110110111101","0000111000101110001011100010","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000110110011101100111011001","0000110111001101110011011100","0000110101011101010111010101","0000110000101100001011000010","0000110000011100000111000001","0000100101011001010110010101","0000100000111000001110000011","0000001100100011001000110010","0000010111100101111001011110","0000100001011000010110000101","0000011101000111010001110100","0000001011110010111100101111","0000001010000010100000101000","0000100000111000001110000011","0000100010101000101010001010","0000011110000111100001111000","0000101101011011010110110101","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111010101110101011101010","0000110110111101101111011011","0000110000101100001011000010","0000110100001101000011010000","0001000000000000000000000000","0000010101100101011001010110","0001000000000000000000000000","0000100101111001011110010111","0000000001110000011100000111","0000001000010010000100100001","0000100010101000101010001010","0000110001111100011111000111","0000101111011011110110111101","0000101111111011111110111111","0000111111001111110011111100","0000111100111111001111110011","0000101010111010101110101011","0000101010101010101010101010","0000110010111100101111001011","0000110011011100110111001101","0000101111001011110010111100","0000111000111110001111100011","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111100001111000011110000","0000111000001110000011100000","0000111000111110001111100011","0000111001111110011111100111","0000111011101110111011101110","0000111101001111010011110100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111101001111010011110100","0000111101001111010011110100","0000111000001110000011100000","0000110000001100000011000000","0000111001001110010011100100","0000100011111000111110001111","0000011101110111011101110111","0000011111000111110001111100","0000111000111110001111100011","0000110011001100110011001100","0000011101010111010101110101","0000111000011110000111100001","0000111101001111010011110100","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111100011111000111110001","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000110010011100100111001001","0000100011001000110010001100","0000011001100110011001100110","0000011010100110101001101010","0000101111001011110010111100","0000111110111111101111111011","0000111010111110101111101011","0000111000101110001011100010","0000111110001111100011111000","0000000001010000010100000101","0000001010100010101000101010","0000111111111111111111111111","0000111011001110110011101100","0000111001011110010111100101","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000110101111101011111010111","0000111111101111111011111110","0000111111001111110011111100","0000111001011110010111100101","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000101001101010011010100110","0000010101000101010001010100","0000100011101000111010001110","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000101110111011101110111011","0000111001011110010111100101","0000101100001011000010110000","0000000011010000110100001101","0000110010001100100011001000","0000111111111111111111111111",
		"0000100100001001000010010000","0000101000101010001010100010","0000101011111010111110101111","0000100001001000010010000100","0000100000111000001110000011","0000010010100100101001001010","0000001110100011101000111010","0000101010001010100010101000","0000111000101110001011100010","0000110000101100001011000010","0000111010011110100111101001","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111101001111010011110100","0000111011001110110011101100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111100101111001011110010","0000111101011111010111110101","0000111110111111101111111011","0000100110111001101110011011","0000010000010100000101000001","0000001111110011111100111111","0000011111110111111101111111","0000100110111001101110011011","0000100001011000010110000101","0000011111000111110001111100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111011011110110111101101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111101001111010011110100","0000111001011110010111100101","0000110101111101011111010111","0000110101101101011011010110","0000110100111101001111010011","0000110001011100010111000101","0000111100011111000111110001","0000111100101111001011110010","0000111101011111010111110101","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111101111111011111110111","0000111101011111010111110101","0000111101001111010011110100","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111101001111010011110100","0000111111111111111111111111","0000111100011111000111110001","0000111101101111011011110110","0000110001111100011111000111","0000101000111010001110100011","0000100011011000110110001101","0000100110011001100110011001","0000011101010111010101110101","0000110011011100110111001101","0000011100110111001101110011","0000001001000010010000100100","0000101000111010001110100011","0000011111100111111001111110","0000010100110101001101010011","0000110110111101101111011011","0000111111111111111111111111","0000111101101111011011110110","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000110001101100011011000110","0000110110101101101011011010","0000110110011101100111011001","0000111001101110011011100110","0000000001110000011100000111","0000010010110100101101001011","0000000100110001001100010011","0000011010100110101001101010","0000001110110011101100111011","0000000111000001110000011100","0000011110110111101101111011","0000110000111100001111000011","0000110110001101100011011000","0000100011111000111110001111","0000111010011110100111101001","0000101000001010000010100000","0000101010001010100010101000","0000110000111100001111000011","0000101010001010100010101000","0000110101001101010011010100","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000100010111000101110001011","0000101100001011000010110000","0000111111111111111111111111","0000110100101101001011010010","0000111111111111111111111111","0000111011001110110011101100","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111011011110110111101101","0000100101011001010110010101","0000111010101110101011101010","0000100000111000001110000011","0000110001011100010111000101","0000010100110101001101010011","0000101101011011010110110101","0000110011001100110011001100","0000110000001100000011000000","0000100110111001101110011011","0000111001111110011111100111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111010111110101111101011","0000111111111111111111111111","0000111111001111110011111100","0000101000111010001110100011","0000100010011000100110001001","0000100001011000010110000101","0000011011100110111001101110","0000101100111011001110110011","0000101111101011111010111110","0000110000111100001111000011","0000111000001110000011100000","0000100001011000010110000101","0000000011110000111100001111","0000010100110101001101010011","0000011111110111111101111111","0000011111110111111101111111","0000011111010111110101111101","0000101100001011000010110000","0000101110001011100010111000","0000111000001110000011100000","0000110001101100011011000110","0000111011111110111111101111","0000111011011110110111101101","0000110010111100101111001011","0000111101011111010111110101","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000110000001100000011000000","0000011000100110001001100010","0000001111100011111000111110","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101101001011010010110100","0000111110111111101111111011","0000001100010011000100110001","0000001101110011011100110111","0000111111001111110011111100","0000111111001111110011111100",
		"0000101001111010011110100111","0000100101111001011110010111","0000100101101001011010010110","0000100000001000000010000000","0000011110110111101101111011","0000010011100100111001001110","0001000000000000000000000000","0000110101101101011011010110","0000110110011101100111011001","0000110010011100100111001001","0000110011011100110111001101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111011111110111111101111","0000111101011111010111110101","0000111101001111010011110100","0000111101001111010011110100","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100011111000111110001","0000101010101010101010101010","0000100100001001000010010000","0000000001000000010000000100","0000001011000010110000101100","0000100001101000011010000110","0000011110100111101001111010","0000101101101011011010110110","0000101110001011100010111000","0000111011001110110011101100","0000111000011110000111100001","0000110011101100111011001110","0000111110011111100111111001","0000111011011110110111101101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111011111110111111101111","0000111011111110111111101111","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111101011111010111110101","0000111101001111010011110100","0000111101011111010111110101","0000111101111111011111110111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111110101111101011111010","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000110110111101101111011011","0000101101001011010010110100","0000101100001011000010110000","0000110011111100111111001111","0000111000001110000011100000","0000110111101101111011011110","0000100111101001111010011110","0000001000100010001000100010","0000001011110010111100101111","0000010101100101011001010110","0000100110011001100110011001","0000110100101101001011010010","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111100101111001011110010","0000110101101101011011010110","0000101111101011111010111110","0000101111101011111010111110","0000110010101100101011001010","0000001001100010011000100110","0000001110000011100000111000","0001000000000000000000000000","0000001010110010101100101011","0000010101000101010001010100","0000001101000011010000110100","0000010001000100010001000100","0000111011101110111011101110","0000110110101101101011011010","0000101110011011100110111001","0000011100000111000001110000","0000011101110111011101110111","0000100100001001000010010000","0000101110001011100010111000","0000101111101011111010111110","0000111000011110000111100001","0000111101001111010011110100","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000110111001101110011011100","0000100110011001100110011001","0000101101111011011110110111","0000111011101110111011101110","0000110110001101100011011000","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111101101111011011110110","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111000001110000011100000","0000110100001101000011010000","0000110100001101000011010000","0000110110111101101111011011","0000101110011011100110111001","0000101100001011000010110000","0001000000000000000000000000","0000110111001101110011011100","0000110001111100011111000111","0000011111010111110101111101","0000101001101010011010100110","0000111111011111110111111101","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000111011111110111111101111","0000111110101111101011111010","0000101111111011111110111111","0000101100011011000110110001","0000011100110111001101110011","0000011111100111111001111110","0000110001111100011111000111","0000011111000111110001111100","0000010110110101101101011011","0000011111100111111001111110","0000100101011001010110010101","0000000010110000101100001011","0000011000100110001001100010","0000010010100100101001001010","0000100000011000000110000001","0000011001010110010101100101","0000011100000111000001110000","0000100011111000111110001111","0000100101011001010110010101","0000011111100111111001111110","0000100000001000000010000000","0000100010011000100110001001","0000111001101110011011100110","0000101011001010110010101100","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000101001001010010010100100","0001000000000000000000000000","0000011111000111110001111100","0000101011011010110110101101","0000111011101110111011101110","0000111111111111111111111111","0000101110101011101010111010","0000101001101010011010100110","0000001100100011001000110010","0000001110110011101100111011","0000111111001111110011111100","0000111111001111110011111100",
		"0000110100101101001011010010","0000001101000011010000110100","0000011111000111110001111100","0000100010001000100010001000","0000011011100110111001101110","0000010100000101000001010000","0001000000000000000000000000","0000100101011001010110010101","0000110111111101111111011111","0000110100001101000011010000","0000110010111100101111001011","0000111001101110011011100110","0000111111111111111111111111","0000111100001111000011110000","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000110111111101111111011111","0000100111101001111010011110","0000010011000100110001001100","0000000101000001010000010100","0000010100000101000001010000","0000100010011000100110001001","0000011100100111001001110010","0000101001011010010110100101","0000111000111110001111100011","0000101100111011001110110011","0000100100111001001110010011","0000110100111101001111010011","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111010001110100011101000","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000101111111011111110111111","0000111011111110111111101111","0000110100111101001111010011","0000111010001110100011101000","0000110101011101010111010101","0000111100001111000011110000","0000011110010111100101111001","0000000101010001010100010101","0000011111110111111101111111","0000100011111000111110001111","0000111001011110010111100101","0000111100001111000011110000","0000111101011111010111110101","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000110100001101000011010000","0000111010011110100111101001","0000110010111100101111001011","0000001111100011111000111110","0000000110010001100100011001","0000000010000000100000001000","0000000010110000101100001011","0000001100010011000100110001","0000001000010010000100100001","0000001100010011000100110001","0000100000001000000010000000","0000101100001011000010110000","0000101111111011111110111111","0000010100010101000101010001","0000010111000101110001011100","0000101100011011000110110001","0000000011100000111000001110","0000110011011100110111001101","0000111011101110111011101110","0000111111001111110011111100","0000111111111111111111111111","0000111110011111100111111001","0000111100111111001111110011","0000111101111111011111110111","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111011101110111011101110","0000110101001101010011010100","0000101100011011000110110001","0000111001011110010111100101","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111110001111100011111000","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110111111101111111011","0000111101011111010111110101","0000110100101101001011010010","0000101111101011111010111110","0000110110011101100111011001","0000110000011100000111000001","0000111010111110101111101011","0000011111110111111101111111","0000100010111000101110001011","0000110000111100001111000011","0000101110011011100110111001","0000011010000110100001101000","0000111011011110110111101101","0000111111111111111111111111","0000111110101111101011111010","0000111011011110110111101101","0000111111111111111111111111","0000111100001111000011110000","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111100101111001011110010","0000111101001111010011110100","0000101100001011000010110000","0000011101110111011101110111","0000100000111000001110000011","0000100111011001110110011101","0000111000111110001111100011","0000001110110011101100111011","0000011011000110110001101100","0000010001010100010101000101","0000000100000001000000010000","0000000111110001111100011111","0001000000000000000000000000","0000000011010000110100001101","0000001000000010000000100000","0000001011010010110100101101","0000001010110010101100101011","0000000000110000001100000011","0000001011010010110100101101","0000010001110100011101000111","0000010001100100011001000110","0000010011000100110001001100","0000011010010110100101101001","0000100011001000110010001100","0000111100111111001111110011","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100101111001011110010","0000111001011110010111100101","0000111100001111000011110000","0000111111101111111011111110","0000111010101110101011101010","0000100010111000101110001011","0001000000000000000000000000","0000010000100100001001000010","0000100011011000110110001101","0000101101001011010010110100","0000001101000011010000110100","0000000000100000001000000010","0000000011100000111000001110","0000101000111010001110100011","0000111111001111110011111100","0000111111001111110011111100",
		"0000111101111111011111110111","0001000000000000000000000000","0000011100010111000101110001","0000100000111000001110000011","0000011100010111000101110001","0000010010000100100001001000","0000010000010100000101000001","0000001111100011111000111110","0000110100011101000111010001","0000110011001100110011001100","0000101001111010011110100111","0000100110111001101110011011","0000111001011110010111100101","0000111110111111101111111011","0000111111111111111111111111","0000111100011111000111110001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000101001011010010110100101","0000110110011101100111011001","0000000100010001000100010001","0000000011000000110000001100","0000100100101001001010010010","0000100100011001000110010001","0000100001011000010110000101","0000101011101010111010101110","0000101001001010010010100100","0000011001000110010001100100","0000101010101010101010101010","0000110011111100111111001111","0000111110101111101011111010","0000111100011111000111110001","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111110011111100111111001","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111110101111101011111010","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111001001110010011100100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000111110011111100111111001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000110000011100000111000001","0000111101001111010011110100","0000110110001101100011011000","0000111000101110001011100010","0000111000111110001111100011","0000111001111110011111100111","0000110110001101100011011000","0000100011001000110010001100","0000001110100011101000111010","0000011101010111010101110101","0000101111111011111110111111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000110011101100111011001110","0000111111101111111011111110","0000111111111111111111111111","0000010111000101110001011100","0001000000000000000000000000","0000000001000000010000000100","0000000101100001011000010110","0000000000010000000100000001","0000000011100000111000001110","0000010001110100011101000111","0000010110000101100001011000","0000011101110111011101110111","0000010010110100101101001011","0000010110100101101001011010","0000001111100011111000111110","0000000101100001011000010110","0000010101010101010101010101","0000111000001110000011100000","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000110011111100111111001111","0000101100001011000010110000","0000011001010110010101100101","0000110001001100010011000100","0000111010011110100111101001","0000111010011110100111101001","0000111010011110100111101001","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110101011101010111010101","0000101110101011101010111010","0000110011001100110011001100","0000110111001101110011011100","0000110111101101111011011110","0000111011001110110011101100","0000000001010000010100000101","0000011111110111111101111111","0000110100101101001011010010","0000100100011001000110010001","0000100110001001100010011000","0000111110001111100011111000","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110011111100111111001","0000110011101100111011001110","0000101111001011110010111100","0000100011001000110010001100","0000011000100110001001100010","0000101000001010000010100000","0000100100101001001010010010","0000011101100111011001110110","0000011010010110100101101001","0000001100010011000100110001","0000001101110011011100110111","0000011010110110101101101011","0000010111010101110101011101","0000011100110111001101110011","0000011001100110011001100110","0000100000101000001010000010","0000011000010110000101100001","0000100000001000000010000000","0000100011011000110110001101","0000010011110100111101001111","0000000101110001011100010111","0000000010000000100000001000","0000001101010011010100110101","0000010110100101101001011010","0000011000100110001001100010","0000101110011011100110111001","0000110011111100111111001111","0000110011111100111111001111","0000110110001101100011011000","0000101010111010101110101011","0000101110111011101110111011","0000110101001101010011010100","0000111111011111110111111101","0000111110011111100111111001","0000110111111101111111011111","0000100100001001000010010000","0000010010100100101001001010","0000000010110000101100001011","0001000000000000000000000000","0000010011010100110101001101","0000000110010001100100011001","0000000011000000110000001100","0000100010011000100110001001","0000111111011111110111111101","0000111111011111110111111101",
		"0000111111111111111111111111","0000010010110100101101001011","0000010101100101011001010110","0000011110110111101101111011","0000100000101000001010000010","0000010010010100100101001001","0000011001100110011001100110","0000010010000100100001001000","0000001110100011101000111010","0000100110011001100110011001","0000100101111001011110010111","0000100011101000111010001110","0000100011011000110110001101","0000110010101100101011001010","0000111100001111000011110000","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111101111111011111110111","0000111110101111101011111010","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111110101111101011111010","0000111010011110100111101001","0000110101001101010011010100","0000100010101000101010001010","0001000000000000000000000000","0000001100110011001100110011","0000101100001011000010110000","0000101000101010001010100010","0000100010101000101010001010","0000011101010111010101110101","0000011111110111111101111111","0000011110010111100101111001","0000100001101000011010000110","0000100101011001010110010101","0000111011111110111111101111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111110111111101111111011","0000111110101111101011111010","0000111110011111100111111001","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000110111111101111111011111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000110100111101001111010011","0000111111111111111111111111","0000111000101110001011100010","0000111111011111110111111101","0000111101101111011011110110","0000111010111110101111101011","0000111111111111111111111111","0000110101101101011011010110","0000110011001100110011001100","0000001010100010101000101010","0000101001001010010010100100","0000110101111101011111010111","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111100101111001011110010","0000110010001100100011001000","0000111101001111010011110100","0000111001111110011111100111","0000011011010110110101101101","0000000000110000001100000011","0000000011100000111000001110","0000011010010110100101101001","0000001011110010111100101111","0000000101100001011000010110","0000000110000001100000011000","0000011010000110100001101000","0000100011001000110010001100","0000001110010011100100111001","0000010100000101000001010000","0000010011110100111101001111","0001000000000000000000000000","0000110001011100010111000101","0000111001111110011111100111","0000111010011110100111101001","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000110111111101111111011111","0000010000000100000001000000","0000000000100000001000000010","0000100000011000000110000001","0000110100001101000011010000","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000101100111011001110110011","0000101111011011110110111101","0000110011111100111111001111","0000011101100111011001110110","0000110111001101110011011100","0000111111111111111111111111","0000011010000110100001101000","0000001000110010001100100011","0000101001001010010010100100","0000100100101001001010010010","0000110010101100101011001010","0000110100011101000111010001","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000100110011001100110011001","0000100111011001110110011101","0000011101100111011001110110","0000011110000111100001111000","0000100101001001010010010100","0000011010000110100001101000","0000010010000100100001001000","0000001100010011000100110001","0000000100000001000000010000","0000011111110111111101111111","0000100110111001101110011011","0000101111001011110010111100","0000101110111011101110111011","0000110011011100110111001101","0000111100111111001111110011","0000111110011111100111111001","0000111001101110011011100110","0000111111111111111111111111","0000111110101111101011111010","0000111000011110000111100001","0000100001111000011110000111","0000001010110010101100101011","0000000110100001101000011010","0000010100000101000001010000","0000010111010101110101011101","0000101010111010101110101011","0000101111011011110110111101","0000101111101011111010111110","0000111011111110111111101111","0000111000101110001011100010","0000111110001111100011111000","0000101110001011100010111000","0000111110111111101111111011","0000111111111111111111111111","0000110100111101001111010011","0000111001101110011011100110","0000110110101101101011011010","0000111100101111001011110010","0000110010001100100011001000","0000011001010110010101100101","0000000100000001000000010000","0000110101011101010111010101","0000111111011111110111111101","0000111111011111110111111101",
		"0000111111001111110011111100","0000101000111010001110100011","0000000111110001111100011111","0000100100101001001010010010","0000100000111000001110000011","0000011000110110001101100011","0000011000100110001001100010","0000010110110101101101011011","0001000000000000000000000000","0000001010100010101000101010","0000010101010101010101010101","0000011110000111100001111000","0000011111010111110101111101","0000100010001000100010001000","0000101100101011001010110010","0000111000011110000111100001","0000111011011110110111101101","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000110001101100011011000110","0000111011101110111011101110","0000011011010110110101101101","0001000000000000000000000000","0000000111110001111100011111","0000110001101100011011000110","0000101111101011111010111110","0000001111110011111100111111","0000011100100111001001110010","0000100010111000101110001011","0000011101110111011101110111","0000010110010101100101011001","0000101011011010110110101101","0000100111011001110110011101","0000101101101011011010110110","0000111110001111100011111000","0000111111111111111111111111","0000111011111110111111101111","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110111111101111111011","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111010101110101011101010","0000111000111110001111100011","0000111110001111100011111000","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111000011110000111100001","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111010001110100011101000","0000111000101110001011100010","0000111010111110101111101011","0000110001101100011011000110","0000111100111111001111110011","0000101010011010100110101001","0000101000011010000110100001","0000110001011100010111000101","0000110111101101111011011110","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111001111110011111100","0000110010111100101111001011","0000100000111000001110000011","0000000100100001001000010010","0001000000000000000000000000","0000010111000101110001011100","0000010010100100101001001010","0000001111100011111000111110","0000010000010100000101000001","0000000011010000110100001101","0000000001010000010100000101","0000000111110001111100011111","0000000000010000000100000001","0000010101000101010001010100","0000111101111111011111110111","0000111001111110011111100111","0000100110111001101110011011","0000111010111110101111101011","0000111101101111011011110110","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111000101110001011100010","0001000000000000000000000000","0000010100110101001101010011","0000110000111100001111000011","0000110011101100111011001110","0000111101101111011011110110","0000110010101100101011001010","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000110110101101101011011010","0000101111001011110010111100","0000101010101010101010101010","0000101000111010001110100011","0000101101011011010110110101","0000101110111011101110111011","0000111100111111001111110011","0000011111000111110001111100","0000000101000001010000010100","0000011011110110111101101111","0000001000000010000000100000","0000110110001101100011011000","0000111001101110011011100110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101011111010111110101","0000111101011111010111110101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111101101111011011110110","0000111010101110101011101010","0000100111001001110010011100","0000101110111011101110111011","0000011111110111111101111111","0000011001100110011001100110","0000010011010100110101001101","0000010010010100100101001001","0000001010100010101000101010","0000001101010011010100110101","0000000001100000011000000110","0000010000100100001001000010","0000100110011001100110011001","0000110101101101011011010110","0000110011101100111011001110","0000101011111010111110101111","0000111011111110111111101111","0000111001011110010111100101","0000110000101100001011000010","0000110010001100100011001000","0000110110101101101011011010","0000111100101111001011110010","0000111111111111111111111111","0000111011101110111011101110","0000111101001111010011110100","0000011000000110000001100000","0001000000000000000000000000","0000010000000100000001000000","0000101000001010000010100000","0000110000001100000011000000","0000110001001100010011000100","0000110000111100001111000011","0000111001001110010011100100","0000111111111111111111111111","0000110101011101010111010101","0000110010011100100111001001","0000111010101110101011101010","0000110111101101111011011110","0000110001101100011011000110","0000111111111111111111111111","0000111111111111111111111111","0000101010101010101010101010","0000001000110010001100100011","0000001000010010000100100001","0000111001011110010111100101","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111111111111111111111","0000110100101101001011010010","0000000110010001100100011001","0000100101111001011110010111","0000011100010111000101110001","0000011011100110111001101110","0000011001100110011001100110","0000011100010111000101110001","0000010111000101110001011100","0000000100000001000000010000","0000000011110000111100001111","0000001011110010111100101111","0000011110100111101001111010","0000100000101000001010000010","0000100011111000111110001111","0000100011101000111010001110","0000101010011010100110101001","0000110001111100011111000111","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000110010101100101011001010","0000111111111111111111111111","0000011101000111010001110100","0000000001000000010000000100","0000010111100101111001011110","0000110100111101001111010011","0000010111000101110001011100","0000010010100100101001001010","0000101100001011000010110000","0000010111000101110001011100","0000100100001001000010010000","0000011001100110011001100110","0000010101000101010001010100","0000011101010111010101110101","0000110001011100010111000101","0000110110101101101011011010","0000110001011100010111000101","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111110111111101111111011","0000111110101111101011111010","0000111110001111100011111000","0000111101111111011111110111","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111100101111001011110010","0000110100101101001011010010","0000111010111110101111101011","0000111101011111010111110101","0000111101101111011011110110","0000111110111111101111111011","0000111011111110111111101111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000110111001101110011011100","0000110111001101110011011100","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000110111001101110011011100","0000111110111111101111111011","0000111101111111011111110111","0000111101111111011111110111","0000111111111111111111111111","0000110010111100101111001011","0000110110111101101111011011","0000101111111011111110111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000100101011001010110010101","0000011110010111100101111001","0000000111110001111100011111","0000000011000000110000001100","0000010000010100000101000001","0000010101100101011001010110","0000001111110011111100111111","0000010111000101110001011100","0000101101111011011110110111","0000011100000111000001110000","0000011101000111010001110100","0000011011100110111001101110","0000110101011101010111010101","0000101001001010010010100100","0000011101000111010001110100","0000111011111110111111101111","0000111110001111100011111000","0000111111011111110111111101","0000111111101111111011111110","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111010111110101111101011","0000000010110000101100001011","0000000111110001111100011111","0000100000101000001010000010","0000111101011111010111110101","0000111011001110110011101100","0000101100011011000110110001","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111111101111111011111110","0000111011111110111111101111","0000110011111100111111001111","0000101010001010100010101000","0000100011001000110010001100","0000100000101000001010000010","0000100011011000110110001101","0000100011111000111110001111","0000110010011100100111001001","0000011000010110000101100001","0001000000000000000000000000","0000010101100101011001010110","0000000000100000001000000010","0000111000101110001011100010","0000111100011111000111110001","0000111101001111010011110100","0000111100001111000011110000","0000111111101111111011111110","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111111111111111111111111","0000100000001000000010000000","0000110001111100011111000111","0000110001111100011111000111","0000101100001011000010110000","0000101101001011010010110100","0000111010001110100011101000","0000101010011010100110101001","0000010100010101000101010001","0001000000000000000000000000","0000001110110011101100111011","0000100011111000111110001111","0000101110101011101010111010","0000111011111110111111101111","0000110011101100111011001110","0000111111111111111111111111","0000110100111101001111010011","0000101001111010011110100111","0000101110011011100110111001","0000110100001101000011010000","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111100001111000011110000","0000110010011100100111001001","0000011100100111001001110010","0000010100000101000001010000","0000010111010101110101011101","0000100010011000100110001001","0000110011111100111111001111","0000110110101101101011011010","0000101101111011011110110111","0000111010011110100111101001","0000111101011111010111110101","0000110111111101111111011111","0000111000111110001111100011","0000110110101101101011011010","0000101110001011100010111000","0000111000001110000011100000","0000111110001111100011111000","0000011011110110111101101111","0000001000100010001000100010","0000010100110101001101010011","0000111100101111001011110010","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111111111111111111111","0000111111111111111111111111","0000010010010100100101001001","0000011101000111010001110100","0000011000110110001101100011","0000010111010101110101011101","0000011100100111001001110010","0000101100101011001010110010","0000011101100111011001110110","0000011110000111100001111000","0000011011110110111101101111","0000001101000011010000110100","0001000000000000000000000000","0000001111000011110000111100","0000011110010111100101111001","0000101001101010011010100110","0000101000001010000010100000","0000100111101001111010011110","0000101000001010000010100000","0000101010011010100110101001","0000101111001011110010111100","0000110101011101010111010101","0000111011011110110111101101","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111001101110011011100110","0000011111100111111001111110","0000000010110000101100001011","0000100111011001110110011101","0000100010101000101010001010","0000100001111000011110000111","0000011010000110100001101000","0000010100000101000001010000","0000101000011010000110100001","0000100010001000100010001000","0000011011110110111101101111","0000101001011010010110100101","0000101000011010000110100001","0000100011111000111110001111","0000101011001010110010101100","0000111011101110111011101110","0000111110111111101111111011","0000111011011110110111101101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111101111111011111110111","0000111101011111010111110101","0000111100111111001111110011","0000111100101111001011110010","0000111100111111001111110011","0000111111111111111111111111","0000111011101110111011101110","0000110000101100001011000010","0000111100011111000111110001","0000111100111111001111110011","0000111100101111001011110010","0000111110001111100011111000","0000111110101111101011111010","0000111111011111110111111101","0000111110011111100111111001","0000111001011110010111100101","0000111111111111111111111111","0000111101111111011111110111","0000110111101101111011011110","0000101101101011011010110110","0000111100001111000011110000","0000111101111111011111110111","0000111100101111001011110010","0000101110011011100110111001","0000111111001111110011111100","0000111010111110101111101011","0000111111101111111011111110","0000111101001111010011110100","0000110111101101111011011110","0000111001111110011111100111","0000101001101010011010100110","0000111111111111111111111111","0000111011111110111111101111","0000111101011111010111110101","0000111110111111101111111011","0000111100001111000011110000","0000100000011000000110000001","0000011100000111000001110000","0000000101010001010100010101","0000000110110001101100011011","0000001000100010001000100010","0000011010100110101001101010","0000001110000011100000111000","0000010101010101010101010101","0000011100000111000001110000","0000011010100110101001101010","0000011010010110100101101001","0000011010010110100101101001","0000100110001001100010011000","0000100001011000010110000101","0000110111111101111111011111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000100000101000001010000010","0000000001100000011000000110","0000001001010010010100100101","0000100101011001010110010101","0000111110001111100011111000","0000101010111010101110101011","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000101101001011010010110100","0000100100101001001010010010","0000100010111000101110001011","0000100100011001000110010001","0000100010001000100010001000","0000010101000101010001010100","0000101101001011010010110100","0000010110010101100101011001","0000000011010000110100001101","0000010000000100000001000000","0000000110000001100000011000","0000110101001101010011010100","0000111101111111011111110111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111100101111001011110010","0000111100001111000011110000","0000111101001111010011110100","0000111111111111111111111111","0000101010001010100010101000","0000110000011100000111000001","0000111110001111100011111000","0000110101001101010011010100","0000111000001110000011100000","0000111010101110101011101010","0000101101101011011010110110","0000011011000110110001101100","0000001101100011011000110110","0000000101100001011000010110","0000011001110110011101100111","0000100000011000000110000001","0000101000001010000010100000","0000100110001001100010011000","0000100011101000111010001110","0000010000110100001101000011","0000010110000101100001011000","0000101110011011100110111001","0000111010111110101111101011","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000110101101101011011010110","0000101100011011000110110001","0000010101110101011101010111","0000100110011001100110011001","0000100111011001110110011101","0000100110001001100010011000","0000101010101010101010101010","0000100110111001101110011011","0000111100101111001011110010","0000111001101110011011100110","0000111000011110000111100001","0000101111111011111110111111","0000101011101010111010101110","0000110110001101100011011000","0000110110011101100111011001","0000011111110111111101111111","0000001111010011110100111101","0000100110101001101010011010","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110",
		"0000111111011111110111111101","0000111101111111011111110111","0000101011011010110110101101","0000001110100011101000111010","0000100001101000011010000110","0000010111100101111001011110","0000001111010011110100111101","0000011000110110001101100011","0000011110110111101101111011","0000101100011011000110110001","0000101000001010000010100000","0000110010101100101011001010","0000101000101010001010100010","0001000000000000000000000000","0001000000000000000000000000","0000100010101000101010001010","0000100010011000100110001001","0000011110110111101101111011","0000100101011001010110010101","0000110000111100001111000011","0000110111101101111011011110","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000010110110101101101011011","0000010000000100000001000000","0000101101001011010010110100","0000010001010100010101000101","0000011001100110011001100110","0000100101101001011010010110","0000101101001011010010110100","0000010001110100011101000111","0000011101110111011101110111","0000110001001100010011000100","0000100111011001110110011101","0000011110000111100001111000","0000110010011100100111001001","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000111101111111011111110111","0000111010011110100111101001","0000111101001111010011110100","0000111001101110011011100110","0000111001101110011011100110","0000110110111101101111011011","0000110100011101000111010001","0000110101011101010111010101","0000101100101011001010110010","0000101111001011110010111100","0000110001101100011011000110","0000111010011110100111101001","0000111101001111010011110100","0000101111011011110110111101","0000111100111111001111110011","0000110000011100000111000001","0000111111111111111111111111","0000111110001111100011111000","0000101101011011010110110101","0000100111101001111010011110","0000110100001101000011010000","0000111001111110011111100111","0000101101001011010010110100","0000101100011011000110110001","0000111100011111000111110001","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000101011011010110110101101","0000111010001110100011101000","0000111100001111000011110000","0000111001111110011111100111","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111100101111001011110010","0000111101111111011111110111","0000100111001001110010011100","0000111100101111001011110010","0000111100001111000011110000","0000111110111111101111111011","0000111111111111111111111111","0000111001111110011111100111","0000011100010111000101110001","0000011010100110101001101010","0000000011010000110100001101","0000000001110000011100000111","0000011001100110011001100110","0000110000101100001011000010","0000001000110010001100100011","0000011011110110111101101111","0000011010100110101001101010","0000100000011000000110000001","0000011011110110111101101111","0000101001111010011110100111","0000100011101000111010001110","0000101000111010001110100011","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000001001100010011000100110","0000000110010001100100011001","0000001100000011000000110000","0000111010111110101111101011","0000101111101011111010111110","0000101001111010011110100111","0000110010001100100011001000","0000111000111110001111100011","0000110100011101000111010001","0000101011111010111110101111","0000110000111100001111000011","0000101110001011100010111000","0000101010001010100010101000","0000011110000111100001111000","0000011001100110011001100110","0000011100100111001001110010","0000011110100111101001111010","0000010011100100111001001110","0000001000000010000000100000","0000010010010100100101001001","0000011101010111010101110101","0000110010001100100011001000","0000111111001111110011111100","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111011111110111111101111","0000111100011111000111110001","0000111111111111111111111111","0000111111011111110111111101","0000110100101101001011010010","0000100011011000110110001101","0000111110001111100011111000","0000110100101101001011010010","0000111011011110110111101101","0000111111001111110011111100","0000110010111100101111001011","0000110111101101111011011110","0000010101000101010001010100","0000000000010000000100000001","0000010010110100101101001011","0000010100110101001101010011","0000010111100101111001011110","0000011000010110000101100001","0000100000101000001010000010","0000010000110100001101000011","0000000111110001111100011111","0000011000110110001101100011","0000100100111001001110010011","0000111000111110001111100011","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111011101110111011101110","0000101110011011100110111001","0000101111111011111110111111","0000110111001101110011011100","0000110111111101111111011111","0000110110111101101111011011","0000111011001110110011101100","0000110111011101110111011101","0000110111111101111111011111","0000101001011010010110100101","0000101100011011000110110001","0000110000111100001111000011","0000110100011101000111010001","0000100010111000101110001011","0001000000000000000000000000","0000111000001110000011100000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111100101111001011110010","0000111011001110110011101100","0000000110100001101000011010","0000100101101001011010010110","0000010001110100011101000111","0000011000000110000001100000","0000001110100011101000111010","0000011110010111100101111001","0000100011111000111110001111","0000100100011001000110010001","0000101000111010001110100011","0000101011101010111010101110","0000101011111010111110101111","0000011111010111110101111101","0000000001110000011100000111","0000000100000001000000010000","0000011110110111101101111011","0000100101001001010010010100","0000011110110111101101111011","0000100111011001110110011101","0000110001111100011111000111","0000111000111110001111100011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111011101110111011101110","0000111010111110101111101011","0000111111111111111111111111","0000111011111110111111101111","0000110111111101111111011111","0000111010001110100011101000","0000001010110010101100101011","0000011000100110001001100010","0000100111111001111110011111","0000001011100010111000101110","0000011100100111001001110010","0000101101001011010010110100","0000100111001001110010011100","0000110001111100011111000111","0000101001001010010010100100","0000011101000111010001110100","0000101111101011111010111110","0000111111111111111111111111","0000111111011111110111111101","0000110110011101100111011001","0000110110001101100011011000","0000101111001011110010111100","0000101101001011010010110100","0000101011101010111010101110","0000100101001001010010010100","0000011111000111110001111100","0000100100011001000110010001","0000101010001010100010101000","0000101111001011110010111100","0000111100001111000011110000","0000111110011111100111111001","0000111101011111010111110101","0000101111101011111010111110","0000101010111010101110101011","0000110000101100001011000010","0000110011101100111011001110","0000110011111100111111001111","0000110010101100101011001010","0000100011101000111010001110","0000100001111000011110000111","0000111001111110011111100111","0000110000101100001011000010","0000011001110110011101100111","0000111000011110000111100001","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111101111111011111110","0000111001101110011011100110","0000110101111101011111010111","0000101000011010000110100001","0000111111111111111111111111","0000111000011110000111100001","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111000001110000011100000","0000101001101010011010100110","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111001011110010111100101","0000111000001110000011100000","0000011101000111010001110100","0000011010010110100101101001","0001000000000000000000000000","0000000011010000110100001101","0000010011110100111101001111","0000101011001010110010101100","0000010111000101110001011100","0000101111001011110010111100","0000101001001010010010100100","0000100110001001100010011000","0000011010010110100101101001","0000011101100111011001110110","0000101011111010111110101111","0000111111101111111011111110","0000111110001111100011111000","0000111110001111100011111000","0000111111111111111111111111","0000111101101111011011110110","0000111000011110000111100001","0000110111111101111111011111","0000111001101110011011100110","0000111000111110001111100011","0000101111001011110010111100","0000100101101001011010010110","0000000101010001010100010101","0000000011110000111100001111","0000000101000001010000010100","0000100101001001010010010100","0000110101111101011111010111","0000100010111000101110001011","0000101100001011000010110000","0000101010101010101010101010","0000110010101100101011001010","0000110110001101100011011000","0000111111111111111111111111","0000110101101101011011010110","0000101000101010001010100010","0000100100111001001110010011","0000010100010101000101010001","0000011010010110100101101001","0000010100010101000101010001","0000011100010111000101110001","0001000000000000000000000000","0000001000100010001000100010","0000011101110111011101110111","0000011010010110100101101001","0000111000101110001011100010","0000111111111111111111111111","0000111111001111110011111100","0000111000001110000011100000","0000111111111111111111111111","0000111110011111100111111001","0000111111011111110111111101","0000111100011111000111110001","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000110101001101010011010100","0000110001011100010111000101","0000111111111111111111111111","0000111000101110001011100010","0000111100101111001011110010","0000111111011111110111111101","0000110011101100111011001110","0000011010110110101101101011","0000010011010100110101001101","0000000010000000100000001000","0000001111000011110000111100","0000010111000101110001011100","0000001000100010001000100010","0000010011100100111001001110","0000001011100010111000101110","0000010100110101001101010011","0000100000001000000010000000","0000100011111000111110001111","0000011101110111011101110111","0000100010011000100110001001","0000100111111001111110011111","0000110100001101000011010000","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111010011110100111101001","0000111001001110010011100100","0000111010111110101111101011","0000111011001110110011101100","0000101010001010100010101000","0000110100011101000111010001","0000110011101100111011001110","0000101110101011101010111010","0000101001111010011110100111","0000100011001000110010001100","0000011000010110000101100001","0000010010110100101101001011","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111111111111111111111111","0000111011001110110011101100","0000011101100111011001110110","0000001100000011000000110000","0000010111010101110101011101","0000001101100011011000110110","0000011111100111111001111110","0000110011001100110011001100","0000011100100111001001110010","0000100011001000110010001100","0000110000101100001011000010","0000101110101011101010111010","0000110011001100110011001100","0000111000001110000011100000","0000101011001010110010101100","0000010000100100001001000010","0001000000000000000000000000","0000000011100000111000001110","0000010110000101100001011000","0000100000011000000110000001","0000101110111011101110111011","0000110111101101111011011110","0000101110101011101010111010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000110111101101111011011110","0000101100101011001010110010","0000111000011110000111100001","0001000000000000000000000000","0000011000100110001001100010","0000100100011001000110010001","0000011001000110010001100100","0000001111110011111100111111","0000010010000100100001001000","0000011101000111010001110100","0000010100100101001001010010","0000010101110101011101010111","0000100100111001001110010011","0000100100011001000110010001","0000100100111001001110010011","0000100011001000110010001100","0000100000001000000010000000","0000011111000111110001111100","0000100101101001011010010110","0000101110111011101110111011","0000110101111101011111010111","0000110100111101001111010011","0000110011101100111011001110","0000110010101100101011001010","0000110101111101011111010111","0000111111111111111111111111","0000111101001111010011110100","0000110001011100010111000101","0000110010101100101011001010","0000011100000111000001110000","0000111000001110000011100000","0000100110101001101010011010","0000100110001001100010011000","0000011011100110111001101110","0000011100000111000001110000","0000110001101100011011000110","0000011001110110011101100111","0000011110000111100001111000","0000111101001111010011110100","0000111111111111111111111111","0000111000111110001111100011","0000110111011101110111011101","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111101101111011011110110","0000111000011110000111100001","0000110101011101010111010101","0000101001101010011010100110","0000111000001110000011100000","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111110101111101011111010","0000111010101110101011101010","0000111111111111111111111111","0000100101001001010010010100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111000001110000011100000","0000101110011011100110111001","0000100001111000011110000111","0000011001100110011001100110","0001000000000000000000000000","0001000000000000000000000000","0000010100100101001001010010","0000011010000110100001101000","0000011101100111011001110110","0000110110001101100011011000","0000110110111101101111011011","0000110100011101000111010001","0000011101010111010101110101","0000010101110101011101010111","0000110111001101110011011100","0000111100001111000011110000","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000111111111111111111111111","0000111011001110110011101100","0000110111011101110111011101","0000110001111100011111000111","0000110011001100110011001100","0000100010011000100110001001","0000010010010100100101001001","0000000001110000011100000111","0000010110000101100001011000","0000011101000111010001110100","0000101001101010011010100110","0000011101110111011101110111","0000110111111101111111011111","0000110101111101011111010111","0000111101101111011011110110","0000111110001111100011111000","0000110111101101111011011110","0000111001001110010011100100","0000101110011011100110111001","0000011101110111011101110111","0000010100100101001001010010","0000010011110100111101001111","0000010000110100001101000011","0000011010100110101001101010","0001000000000000000000000000","0000001100010011000100110001","0000011000110110001101100011","0000100101101001011010010110","0000011100010111000101110001","0000101101111011011110110111","0000110001001100010011000100","0000111010001110100011101000","0000111110111111101111111011","0000111100101111001011110010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111100111111001111110011","0000111111001111110011111100","0000111010011110100111101001","0000111100011111000111110001","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000100110101001101010011010","0000100010001000100010001000","0000010110100101101001011010","0000000000010000000100000001","0000010001000100010001000100","0000000101100001011000010110","0001000000000000000000000000","0000000110110001101100011011","0000001001010010010100100101","0000010111110101111101011111","0000101101011011010110110101","0000110110011101100111011001","0000110001111100011111000111","0000110100001101000011010000","0000100110111001101110011011","0000101101001011010010110100","0000100010101000101010001010","0000101111111011111110111111","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100001101000011010000","0000111001101110011011100110","0000110010101100101011001010","0000101100001011000010110000","0000110010001100100011001000","0000101000101010001010100010","0000011010100110101001101010","0000100010111000101110001011","0001000000000000000000000000","0000100111101001111010011110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000110100001101000011010000","0000000000010000000100000001","0000011000100110001001100010","0000000011000000110000001100","0000110010111100101111001011","0000111110001111100011111000","0000101110101011101010111010","0000110111011101110111011101","0000110101111101011111010111","0000110011101100111011001110","0000111101011111010111110101","0000111111111111111111111111","0000111110101111101011111010","0000111100001111000011110000","0000111111111111111111111111","0000101100111011001110110011","0000010000100100001001000010","0000010010100100101001001010","0000100000111000001110000011","0000100101101001011010010110","0000100111101001111010011110","0000100101111001011110010111","0000111111111111111111111111","0000111111001111110011111100","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000101001111010011110100111","0000110101101101011011010110","0000101100101011001010110010","0001000000000000000000000000","0000010000010100000101000001","0000101011101010111010101110","0000100101111001011110010111","0000011110100111101001111010","0000100111111001111110011111","0000011000100110001001100010","0000100100101001001010010010","0000101101011011010110110101","0000100101111001011110010111","0000010101100101011001010110","0000011001100110011001100110","0000011110100111101001111010","0000100110011001100110011001","0000101101011011010110110101","0000100110001001100010011000","0000010110110101101101011011","0000001000110010001100100011","0000000010110000101100001011","0000001110000011100000111000","0000010100100101001001010010","0000000011010000110100001101","0000001001100010011000100110","0000001110100011101000111010","0000001111110011111100111111","0000001000010010000100100001","0000001111110011111100111111","0000010101100101011001010110","0000001101110011011100110111","0000000111000001110000011100","0000011011000110110001101100","0000000010000000100000001000","0000100010101000101010001010","0000111111111111111111111111","0000111010101110101011101010","0000111111001111110011111100","0000110000011100000111000001","0000111101011111010111110101","0000111111001111110011111100","0000111110101111101011111010","0000111111001111110011111100","0000111111101111111011111110","0000111111101111111011111110","0000111111001111110011111100","0000111101001111010011110100","0000111010001110100011101000","0000101110111011101110111011","0000101011001010110010101100","0000110011011100110111001101","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111100101111001011110010","0000111100001111000011110000","0000101010111010101110101011","0000111101001111010011110100","0000111111111111111111111111","0000111001011110010111100101","0000111111111111111111111111","0000100010011000100110001001","0000011100110111001101110011","0000010111100101111001011110","0000000110000001100000011000","0000000011010000110100001101","0001000000000000000000000000","0000011101000111010001110100","0000101000001010000010100000","0000011110000111100001111000","0000101100101011001010110010","0000101010101010101010101010","0000100111011001110110011101","0000100101101001011010010110","0000111110111111101111111011","0000111111111111111111111111","0000110100011101000111010001","0000111110101111101011111010","0000111111001111110011111100","0000111100111111001111110011","0000110100011101000111010001","0000101110011011100110111001","0000100111001001110010011100","0000100001001000010010000100","0000001111110011111100111111","0000000001000000010000000100","0000010010110100101101001011","0000101000111010001110100011","0000010111100101111001011110","0000100100001001000010010000","0000110100101101001011010010","0000101011111010111110101111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110011101100111011001","0000100010111000101110001011","0000011001110110011101100111","0000010000110100001101000011","0000001111100011111000111110","0000000010110000101100001011","0000000001110000011100000111","0000010000010100000101000001","0000010111000101110001011100","0000010110010101100101011001","0000010101000101010001010100","0000010100100101001001010010","0000111100111111001111110011","0000101100111011001110110011","0000110100001101000011010000","0000111100011111000111110001","0000111110111111101111111011","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111111001111110011111100","0000111110101111101011111010","0000111111111111111111111111","0000111100011111000111110001","0000111001001110010011100100","0000100000011000000110000001","0000011010100110101001101010","0000011000010110000101100001","0000000001010000010100000101","0000000101010001010100010101","0000000100110001001100010011","0000000100000001000000010000","0000001111100011111000111110","0000011100100111001001110010","0000101011011010110110101101","0000100101111001011110010111","0000100000011000000110000001","0000100000101000001010000010","0000100100101001001010010010","0000110111011101110111011101","0000111110111111101111111011","0000110011101100111011001110","0000111000011110000111100001","0000101010011010100110101001","0000110100011101000111010001","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000110000101100001011000010","0000110111101101111011011110","0000111001111110011111100111","0000101111111011111110111111","0000101101111011011110110111","0000110100111101001111010011","0000101110001011100010111000","0000100010001000100010001000","0000100100001001000010010000","0000010001110100011101000111","0000100000111000001110000011","0001000000000000000000000000","0000111001111110011111100111","0000111100011111000111110001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000111100011111000111110001","0000010001000100010001000100","0000001111010011110100111101","0000000010000000100000001000","0000101110001011100010111000","0000111110011111100111111001","0000101100101011001010110010","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111100111111001111110011","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000110111011101110111011101","0000101101011011010110110101","0000011100110111001101110011","0000001010110010101100101011","0000011010000110100001101000","0000101011111010111110101111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111001101110011011100110","0000111100001111000011110000","0000101000001010000010100000","0000100001101000011010000110","0000100100001001000010010000","0000100000011000000110000001","0000010000100100001001000010","0001000000000000000000000000","0000010100010101000101010001","0000011010100110101001101010","0000010111010101110101011101","0000100000111000001110000011","0000101000011010000110100001","0000011100000111000001110000","0000011100110111001101110011","0000100000011000000110000001","0000010100010101000101010001","0000000001000000010000000100","0001000000000000000000000000","0001000000000000000000000000","0000000000010000000100000001","0000000100110001001100010011","0000000000010000000100000001","0001000000000000000000000000","0000010001000100010001000100","0000100010001000100010001000","0000100110101001101010011010","0000100000011000000110000001","0000010101010101010101010101","0000000001110000011100000111","0000011111010111110101111101","0000010010110100101101001011","0000001100100011001000110010","0000010011010100110101001101","0000011111010111110101111101","0000101110001011100010111000","0000100010111000101110001011","0000111111011111110111111101","0000111101101111011011110110","0000111111001111110011111100","0000100110011001100110011001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111110001111100011111000","0000111111011111110111111101","0000111110111111101111111011","0000111101101111011011110110","0000111101101111011011110110","0000101000011010000110100001","0000101100111011001110110011","0000101100101011001010110010","0000111101011111010111110101","0000111101111111011111110111","0000111011001110110011101100","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111110001111100011111000","0000101110001011100010111000","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000110011101100111011001110","0000101001101010011010100110","0000011100100111001001110010","0000001001000010010000100100","0000000011000000110000001100","0001000000000000000000000000","0000001010010010100100101001","0000010101010101010101010101","0000011110110111101101111011","0000011001010110010101100101","0000101100001011000010110000","0000101101011011010110110101","0000100111011001110110011101","0000101010001010100010101000","0000111111111111111111111111","0000110101111101011111010111","0000111001001110010011100100","0000111101111111011111110111","0000111100011111000111110001","0000111001001110010011100100","0000111110111111101111111011","0000111110101111101011111010","0000101110001011100010111000","0000010010000100100001001000","0000001111010011110100111101","0000011011100110111001101110","0000101111011011110110111101","0000011010100110101001101010","0000011000100110001001100010","0000101001111010011110100111","0000101010011010100110101001","0000110110101101101011011010","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110000011100000111000001","0000100101111001011110010111","0000001110110011101100111011","0000010010000100100001001000","0000001011000010110000101100","0001000000000000000000000000","0000001100100011001000110010","0000100111011001110110011101","0000100010011000100110001001","0000010011100100111001001110","0000010111010101110101011101","0000101000001010000010100000","0000011011110110111101101111","0000010101110101011101010111","0000111111111111111111111111","0000111110001111100011111000","0000111001101110011011100110","0000111110111111101111111011","0000111111011111110111111101","0000111101101111011011110110","0000111101001111010011110100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000110111001101110011011100","0000111111111111111111111111","0000110110011101100111011001","0000100110001001100010011000","0000011010110110101101101011","0000001000110010001100100011","0000001010000010100000101000","0000010011000100110001001100","0000000011000000110000001100","0000000011110000111100001111","0000001100010011000100110001","0000100001111000011110000111","0000100100101001001010010010","0000011010100110101001101010","0000011000110110001101100011","0000100101001001010010010100","0000011011110110111101101111","0000110010101100101011001010","0000101100111011001110110011","0000101011111010111110101111","0000110101001101010011010100","0000110001001100010011000100","0000111011111110111111101111","0000101101111011011110110111","0000111101101111011011110110","0000111111011111110111111101","0000111110111111101111111011","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000110011001100110011001100","0000011101000111010001110100","0000100111011001110110011101","0000101011101010111010101110","0000101001011010010110100101","0000100100111001001110010011","0000100011111000111110001111","0000010000000100000001000000","0000011011010110110101101101","0000001111010011110100111101","0000011001010110010101100101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101101111011011110110","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000100110011001100110011001","0001000000000000000000000000","0000000001010000010100000101","0000100111101001111010011110","0000110011101100111011001110","0000101010101010101010101010","0000111111111111111111111111","0000111110001111100011111000","0000111010101110101011101010","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111100101111001011110010","0000101111101011111010111110","0000011110000111100001111000","0000100000111000001110000011","0000010010000100100001001000","0000101010111010101110101011","0000111101111111011111110111","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000101010101010101010101010","0000011100000111000001110000","0000100001101000011010000110","0000010110100101101001011010","0000100100011001000110010001","0000010111100101111001011110","0000000111110001111100011111","0000000100010001000100010001","0000001011010010110100101101","0000001000000010000000100000","0000001000100010001000100010","0000001000110010001100100011","0000000010110000101100001011","0001000000000000000000000000","0000000011010000110100001101","0000011100100111001001110010","0000011101110111011101110111","0000011000110110001101100011","0000010101010101010101010101","0000100000111000001110000011","0000011100110111001101110011","0000010000100100001001000010","0001000000000000000000000000","0000000010100000101000001010","0000110000111100001111000011","0000100111011001110110011101","0000011011000110110001101100","0000010100100101001001010010","0000100100101001001010010010","0000100010011000100110001001","0000100011011000110110001101","0000101010001010100010101000","0000100111111001111110011111","0000011101100111011001110110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000110111001101110011011100","0000101011101010111010101110","0000111001111110011111100111","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111011011110110111101101","0000111100001111000011110000","0000111111011111110111111101","0000111110101111101011111010","0000111101001111010011110100","0000111111101111111011111110","0000101000111010001110100011","0000101011101010111010101110","0000011111100111111001111110","0000111111111111111111111111","0000111000011110000111100001","0000111010011110100111101001","0000111011101110111011101110","0000111101011111010111110101","0000111010111110101111101011","0000111111111111111111111111","0000110011001100110011001100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101111101011111010111110","0000101000001010000010100000","0000011011010110110101101101","0000001001100010011000100110","0001000000000000000000000000","0000000111000001110000011100","0000000110100001101000011010","0000011000010110000101100001","0000010101100101011001010110","0000010110010101100101011001","0000100001111000011110000111","0000111011001110110011101100","0000100011111000111110001111","0000110101101101011011010110","0000111111111111111111111111","0000101101011011010110110101","0000111111111111111111111111","0000110010111100101111001011","0000110111101101111011011110","0000111110001111100011111000","0000111000011110000111100001","0000011110110111101101111011","0000011011000110110001101100","0000100010001000100010001000","0000100111101001111010011110","0000011101000111010001110100","0000010011000100110001001100","0000011010000110100001101000","0000100110001001100010011000","0000100110001001100010011000","0000111001011110010111100101","0000111111111111111111111111","0000111110001111100011111000","0000110001011100010111000101","0000101110101011101010111010","0000011011000110110001101100","0000010101000101010001010100","0000001010110010101100101011","0000000011000000110000001100","0000000101110001011100010111","0000010110100101101001011010","0000101100011011000110110001","0000010111100101111001011110","0000011110010111100101111001","0000101000001010000010100000","0000010101000101010001010100","0000010110110101101101011011","0000100001111000011110000111","0000101000001010000010100000","0000101110001011100010111000","0000111111111111111111111111","0000111100011111000111110001","0000110111001101110011011100","0000111111011111110111111101","0000111011001110110011101100","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000110000101100001011000010","0000100111011001110110011101","0000011111110111111101111111","0000001010100010101000101010","0001000000000000000000000000","0000000011110000111100001111","0000001110010011100100111001","0000011111010111110101111101","0000110011011100110111001101","0000101110111011101110111011","0000101001101010011010100110","0000101010011010100110101001","0000101100111011001110110011","0000100100001001000010010000","0000100000001000000010000000","0000110100101101001011010010","0000110000111100001111000011","0000111000101110001011100010","0000111010111110101111101011","0000100101111001011110010111","0000111010011110100111101001","0000111010101110101011101010","0000110010011100100111001001","0000110011001100110011001100","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111101101111011011110110","0000011011110110111101101111","0000001011110010111100101111","0000011011110110111101101111","0000100110111001101110011011","0000011101110111011101110111","0000100010011000100110001001","0000001000000010000000100000","0000000011110000111100001111","0000111000101110001011100010","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101101111011011110110","0000111001101110011011100110","0001000000000000000000000000","0000000001110000011100000111","0000100010111000101110001011","0000110101001101010011010100","0000101011101010111010101110","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111101011111010111110101","0000111111111111111111111111","0000111100111111001111110011","0000111101011111010111110101","0000111111111111111111111111","0000111111011111110111111101","0000111011101110111011101110","0000111110111111101111111011","0000111111111111111111111111","0000111010011110100111101001","0000110110101101101011011010","0000110111111101111111011111","0000101101101011011010110110","0000011001010110010101100101","0000100110111001101110011011","0000110101011101010111010101","0000111101011111010111110101","0000111010111110101111101011","0000110100111101001111010011","0000010111010101110101011101","0000011100010111000101110001","0000010100010101000101010001","0000100011001000110010001100","0000011100100111001001110010","0000010110000101100001011000","0000001111010011110100111101","0000001101010011010100110101","0000000010100000101000001010","0000010010000100100001001000","0000011100000111000001110000","0000011111000111110001111100","0000110010011100100111001001","0000111100111111001111110011","0000110101001101010011010100","0000011111110111111101111111","0000100110101001101010011010","0000110101101101011011010110","0000101000111010001110100011","0000001101100011011000110110","0000010011010100110101001101","0000011100000111000001110000","0000001011010010110100101101","0000000010100000101000001010","0000011010100110101001101010","0000010101010101010101010101","0000011111010111110101111101","0000101100111011001110110011","0000101011001010110010101100","0000110000101100001011000010","0000100100101001001010010010","0000100010111000101110001011","0000110010011100100111001001","0000111111011111110111111101","0000111100111111001111110011","0000111110111111101111111011","0000101111101011111010111110","0000110011011100110111001101","0000111101011111010111110101","0000111111111111111111111111","0000111001111110011111100111","0000111010011110100111101001","0000111000101110001011100010","0000111010111110101111101011","0000111111101111111011111110","0000111101111111011111110111","0000111011011110110111101101","0000111110111111101111111011","0000110011101100111011001110","0000011101100111011001110110","0000100001011000010110000101","0000111010001110100011101000","0000110011011100110111001101","0000111110001111100011111000","0000110000011100000111000001","0000111001111110011111100111","0000111011011110110111101101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000110000101100001011000010","0000111010101110101011101010","0000010110110101101101011011","0000100100011001000110010001","0001000000000000000000000000","0000000110010001100100011001","0000010111110101111101011111","0000000100000001000000010000","0000001001110010011100100111","0000011001000110010001100100","0000010000100100001001000010","0000011100000111000001110000","0000110100101101001011010010","0000100000101000001010000010","0000101111011011110110111101","0000101101011011010110110101","0000111111101111111011111110","0000111101101111011011110110","0000111111111111111111111111","0000111111001111110011111100","0000111111011111110111111101","0000111100011111000111110001","0000110100101101001011010010","0000101110101011101010111010","0000101000101010001010100010","0000100010101000101010001010","0000011100010111000101110001","0000011001010110010101100101","0000100101011001010110010101","0000100101111001011110010111","0000110001011100010111000101","0000101010011010100110101001","0000100110011001100110011001","0000010111100101111001011110","0000001001110010011100100111","0000010111000101110001011100","0000001100010011000100110001","0000000011000000110000001100","0000000110010001100100011001","0000001001100010011000100110","0000011110100111101001111010","0000101010111010101110101011","0000011001010110010101100101","0000010110000101100001011000","0000011111000111110001111100","0000100001111000011110000111","0000010111110101111101011111","0000100011111000111110001111","0000011111100111111001111110","0000100001001000010010000100","0000100101001001010010010100","0000101011101010111010101110","0000101111001011110010111100","0000101111111011111110111111","0000101011101010111010101110","0000111011011110110111101101","0000111001101110011011100110","0000111000101110001011100010","0000110111001101110011011100","0000110101001101010011010100","0000101001111010011110100111","0000011111010111110101111101","0000010110000101100001011000","0000001001010010010100100101","0001000000000000000000000000","0000000111010001110100011101","0000100001101000011010000110","0000110101001101010011010100","0000101010001010100010101000","0000101000011010000110100001","0000101010011010100110101001","0000100110101001101010011010","0000011101010111010101110101","0000100010011000100110001001","0000011110110111101101111011","0000101101101011011010110110","0000101100011011000110110001","0000110001111100011111000111","0000110000011100000111000001","0000101101011011010110110101","0000111100101111001011110010","0000101100011011000110110001","0000111110001111100011111000","0000111011001110110011101100","0000110001001100010011000100","0000111001111110011111100111","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111101001111010011110100","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000110011111100111111001111","0000010111110101111101011111","0000001111110011111100111111","0000011000110110001101100011","0000100010011000100110001001","0000010011100100111001001110","0000011100000111000001110000","0000000111100001111000011110","0000111111111111111111111111","0000111101001111010011110100","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000011001110110011101100111","0001000000000000000000000000","0000011001010110010101100101","0000110000011100000111000001","0000101010101010101010101010","0000111100111111001111110011","0000111100111111001111110011","0000111111111111111111111111","0000111110101111101011111010","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000101110101011101010111010","0000111100101111001011110010","0000100000001000000010000000","0000111011111110111111101111","0000111011011110110111101101","0000111010011110100111101001","0000111111111111111111111111","0000111001111110011111100111","0000100011101000111010001110","0000100001101000011010000110","0000100011001000110010001100","0000100000111000001110000011","0000011101100111011001110110","0000011101100111011001110110","0000100101111001011110010111","0000010010110100101101001011","0000010111010101110101011101","0000101111011011110110111101","0000111000011110000111100001","0000110010101100101011001010","0000110100111101001111010011","0000111011111110111111101111","0000101011101010111010101110","0000100110001001100010011000","0000111000101110001011100010","0000111000001110000011100000","0000100000101000001010000010","0000100111111001111110011111","0000110010011100100111001001","0000100101001001010010010100","0000011101010111010101110101","0000001110000011100000111000","0000000010000000100000001000","0000001110100011101000111010","0000100000001000000010000000","0000100011001000110010001100","0000110000101100001011000010","0000101001011010010110100101","0000110001111100011111000111","0000101000111010001110100011","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100101111001011110010","0000101101001011010010110100","0000110010011100100111001001","0000110111111101111111011111","0000111100001111000011110000","0000110101111101011111010111","0000110111011101110111011101","0000110110111101101111011011","0000111010011110100111101001","0000111111111111111111111111","0000111101001111010011110100","0000111001101110011011100110","0000111101001111010011110100","0000111001001110010011100100","0000011001110110011101100111","0000100010001000100010001000","0000101111101011111010111110","0000111100111111001111110011","0000101110101011101010111010","0000111011011110110111101101","0000101101111011011110110111","0000110100101101001011010010","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111000101110001011100010","0000110101011101010111010101","0000011101110111011101110111","0000011010000110100001101000","0000010010100100101001001010","0000001011100010111000101110","0000001010010010100100101001","0000010011110100111101001111","0000000100110001001100010011","0000001110000011100000111000","0000010010110100101101001011","0000010001100100011001000110","0000011010010110100101101001","0000100110101001101010011010","0000100110001001100010011000","0000011101110111011101110111","0000111001111110011111100111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111001111110011111100111","0000111001101110011011100110","0000101111101011111010111110","0000101000001010000010100000","0000011101010111010101110101","0000011010100110101001101010","0000100110001001100010011000","0000100001101000011010000110","0000100101101001011010010110","0000110001111100011111000111","0000101001111010011110100111","0000100010011000100110001001","0000011011100110111001101110","0000010010010100100101001001","0000000100010001000100010001","0000001100010011000100110001","0000010011000100110001001100","0000010110110101101101011011","0000011100000111000001110000","0000011111100111111001111110","0000010000100100001001000010","0000011100000111000001110000","0000011100100111001001110010","0000011110010111100101111001","0000100000111000001110000011","0000101100101011001010110010","0000011010110110101101101011","0000011111110111111101111111","0000010100100101001001010010","0000010010110100101101001011","0000011011100110111001101110","0000100100101001001010010010","0000100111101001111010011110","0000100101101001011010010110","0000100100011001000110010001","0000101111001011110010111100","0000100110101001101010011010","0000010010000100100001001000","0000001111010011110100111101","0000010100000101000001010000","0000000011000000110000001100","0000000000100000001000000010","0001000000000000000000000000","0000011010100110101001101010","0000101100011011000110110001","0000101100111011001110110011","0000101000011010000110100001","0000100100101001001010010010","0000101010001010100010101000","0000100010011000100110001001","0000100100111001001110010011","0000100110111001101110011011","0000100110111001101110011011","0000101011101010111010101110","0000110001101100011011000110","0000110010001100100011001000","0000110011001100110011001100","0000100101011001010110010101","0000101111101011111010111110","0000110001011100010111000101","0000111111111111111111111111","0000101110111011101110111011","0000111111111111111111111111","0000110110011101100111011001","0000110100111101001111010011","0000111111101111111011111110","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111001111110011111100111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000100000001000000010000000","0000010100100101001001010010","0000001101010011010100110101","0000010111000101110001011100","0000100100001001000010010000","0000011000100110001001100010","0000110000011100000111000001","0000111011111110111111101111","0000111110001111100011111000","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111101111111011111110","0000111111111111111111111111","0000111111001111110011111100","0000111100111111001111110011","0000111111101111111011111110","0000101100001011000010110000","0001000000000000000000000000","0000010101100101011001010110","0000100011001000110010001100","0000100110101001101010011010","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100011111000111110001","0000111110101111101011111010","0000111110111111101111111011","0000110101001101010011010100","0000110011111100111111001111","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000111111001111110011111100","0000110000011100000111000001","0000101111001011110010111100","0000101111111011111110111111","0000111110111111101111111011","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000100011011000110110001101","0000011110110111101101111011","0000101011011010110110101101","0000101001101010011010100110","0000110010111100101111001011","0000110101101101011011010110","0000100011001000110010001100","0000011101100111011001110110","0000110011001100110011001100","0000111010101110101011101010","0000101000011010000110100001","0000110001111100011111000111","0000111111011111110111111101","0000110110001101100011011000","0000101101101011011010110110","0000110100101101001011010010","0000111011101110111011101110","0000100101111001011110010111","0000100111101001111010011110","0000111000111110001111100011","0000111111111111111111111111","0000111010101110101011101010","0000101100111011001110110011","0000101010111010101110101011","0000001100000011000000110000","0001000000000000000000000000","0000100001001000010010000100","0000011000000110000001100000","0000101111101011111010111110","0000110000111100001111000011","0000110001001100010011000100","0000111001001110010011100100","0000111100001111000011110000","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000101101011011010110110101","0000101001001010010010100100","0000110000011100000111000001","0000111010111110101111101011","0000110110101101101011011010","0000111000011110000111100001","0000111011001110110011101100","0000111010011110100111101001","0000111110011111100111111001","0000111100001111000011110000","0000111101001111010011110100","0000110000111100001111000011","0000110010111100101111001011","0000011111000111110001111100","0000010011100100111001001110","0000101110111011101110111011","0000111000001110000011100000","0000101100011011000110110001","0000111101111111011111110111","0000110000011100000111000001","0000101100111011001110110011","0000101010011010100110101001","0000111001101110011011100110","0000111110101111101011111010","0000111100011111000111110001","0000011111110111111101111111","0000011101000111010001110100","0000100100101001001010010010","0000000111100001111000011110","0001000000000000000000000000","0000001111000011110000111100","0000010011010100110101001101","0000001010010010100100101001","0000001101010011010100110101","0000001111000011110000111100","0000010010100100101001001010","0000100011101000111010001110","0000100101011001010110010101","0000101110101011101010111010","0000100011101000111010001110","0000111110101111101011111010","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000110110111101101111011011","0000110001101100011011000110","0000101101101011011010110110","0000100111101001111010011110","0000110011011100110111001101","0000111011011110110111101101","0000111001001110010011100100","0000101100101011001010110010","0000101100101011001010110010","0000001000000010000000100000","0000000010100000101000001010","0000001001100010011000100110","0000001111010011110100111101","0000011001010110010101100101","0000011100000111000001110000","0000011110100111101001111010","0000101110111011101110111011","0000100101111001011110010111","0000100000101000001010000010","0000010111100101111001011110","0000010000010100000101000001","0000110011001100110011001100","0000111100011111000111110001","0000101111101011111010111110","0000011110000111100001111000","0000010011000100110001001100","0000101001111010011110100111","0000101000001010000010100000","0000010011110100111101001111","0000011100100111001001110010","0000100001111000011110000111","0000011100100111001001110010","0000011000110110001101100011","0000010110010101100101011001","0000011110000111100001111000","0000011101100111011001110110","0000011110100111101001111010","0000010110110101101101011011","0000000101110001011100010111","0001000000000000000000000000","0000100100101001001010010010","0000111110101111101011111010","0000110000111100001111000011","0000110001011100010111000101","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000110100101101001011010010","0000110000011100000111000001","0000110101001101010011010100","0000110111001101110011011100","0000101111111011111110111111","0000110100111101001111010011","0000110100011101000111010001","0000111110101111101011111010","0000110001101100011011000110","0000111111011111110111111101","0000110001011100010111000101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110000011100000111000001","0000010111010101110101011101","0000000011110000111100001111","0000010000100100001001000010","0000011111110111111101111111","0000010011010100110101001101","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101111111011111110111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000000100110001001100010011","0000000011100000111000001110","0000011111100111111001111110","0000100010001000100010001000","0000111001001110010011100100","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111111101111111011111110","0000110101111101011111010111","0000101000011010000110100001","0000111111111111111111111111","0000111111011111110111111101","0000111011001110110011101100","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000110110011101100111011001","0000111000111110001111100011","0000100101011001010110010101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000011100100111001001110010","0000011001000110010001100100","0000101101101011011010110110","0000100110101001101010011010","0000110010111100101111001011","0000101001001010010010100100","0000010110100101101001011010","0000110000101100001011000010","0000110111101101111011011110","0000100000001000000010000000","0000111101001111010011110100","0000111111111111111111111111","0000111100101111001011110010","0000110011101100111011001110","0000110000111100001111000011","0000111110111111101111111011","0000101101011011010110110101","0000101010001010100010101000","0000110100011101000111010001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000110100001101000011010000","0000010111010101110101011101","0000000101010001010100010101","0000011000000110000001100000","0000100000001000000010000000","0000100011101000111010001110","0000101110101011101010111010","0000101111101011111010111110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110111111101111111011","0000110111111101111111011111","0000110101101101011011010110","0000100001111000011110000111","0000101001111010011110100111","0000101100101011001010110010","0000110111011101110111011101","0000110011101100111011001110","0000110000001100000011000000","0000110111111101111111011111","0000111111101111111011111110","0000110010101100101011001010","0000111111111111111111111111","0000110011011100110111001101","0000100000111000001110000011","0000011111100111111001111110","0000000101110001011100010111","0000011110000111100001111000","0000111000011110000111100001","0000101010011010100110101001","0000111001001110010011100100","0000111000111110001111100011","0000100110111001101110011011","0000100100011001000110010001","0000011011010110110101101101","0000011010000110100001101000","0000010011110100111101001111","0000100011001000110010001100","0000011111100111111001111110","0000001100100011001000110010","0001000000000000000000000000","0000000100100001001000010010","0000010011000100110001001100","0000001110010011100100111001","0000000001100000011000000110","0000001101110011011100110111","0000001111010011110100111101","0000011010100110101001101010","0000010111110101111101011111","0000100010101000101010001010","0000101100011011000110110001","0000100011001000110010001100","0000111011001110110011101100","0000111010111110101111101011","0000111111111111111111111111","0000111111001111110011111100","0000111011111110111111101111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100101111001011110010","0000110100011101000111010001","0000110110001101100011011000","0000111111111111111111111111","0000111111011111110111111101","0000110100001101000011010000","0000110101101101011011010110","0000011110110111101101111011","0001000000000000000000000000","0000100100001001000010010000","0000110111001101110011011100","0000110111101101111011011110","0000110001001100010011000100","0000111111111111111111111111","0000111011111110111111101111","0000111100111111001111110011","0000100100011001000110010001","0000100010111000101110001011","0000010100010101000101010001","0000100000001000000010000000","0000111101001111010011110100","0000100011101000111010001110","0000100101011001010110010101","0000111001011110010111100101","0000110001101100011011000110","0000011011110110111101101111","0000011001010110010101100101","0000010001100100011001000110","0000100101011001010110010101","0000011011110110111101101111","0000100011101000111010001110","0000011110010111100101111001","0000011111100111111001111110","0000011011100110111001101110","0000011110000111100001111000","0000011001100110011001100110","0000001011000010110000101100","0001000000000000000000000000","0000000100010001000100010001","0000100111101001111010011110","0000111001111110011111100111","0000101100111011001110110011","0000110001001100010011000100","0000111011111110111111101111","0000111101111111011111110111","0000111110101111101011111010","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000111101001111010011110100","0000110010001100100011001000","0000101101111011011110110111","0000111111111111111111111111","0000101111111011111110111111","0000101110001011100010111000","0000110001011100010111000101","0000111100011111000111110001","0000111101101111011011110110","0000111110101111101011111010","0000111011011110110111101101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111011111110111111101","0000111100011111000111110001","0000111111111111111111111111","0000111111001111110011111100","0000110100111101001111010011","0000100111011001110110011101","0000000110110001101100011011","0000000111100001111000011110","0000001111100011111000111110","0000101000111010001110100011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111100111111001111110011","0000111111111111111111111111","0000011010110110101101101011","0001000000000000000000000000","0000011011100110111001101110","0000011110110111101101111011","0000100000111000001110000011","0000110000011100000111000001","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000110011101100111011001110","0000110110011101100111011001","0000111101001111010011110100","0000100101001001010010010100","0000111010001110100011101000","0000111100011111000111110001","0000111101011111010111110101","0000111111111111111111111111","0000111100101111001011110010","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000100011011000110110001101","0000111011111110111111101111","0000111111111111111111111111","0000111111001111110011111100","0000110010111100101111001011","0000011101100111011001110110","0000100000001000000010000000","0000010001000100010001000100","0000100100101001001010010010","0000100101001001010010010100","0000010011010100110101001101","0000011011100110111001101110","0000110101111101011111010111","0000100011001000110010001100","0000111111111111111111111111","0000111101111111011111110111","0000110111111101111111011111","0000111111111111111111111111","0000111110101111101011111010","0000111011001110110011101100","0000111100011111000111110001","0000110100001101000011010000","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111011111110111111101","0000111011011110110111101101","0000010110110101101101011011","0000001111000011110000111100","0000000010010000100100001001","0000100111011001110110011101","0000011111010111110101111101","0000100111011001110110011101","0000110111101101111011011110","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111011101110111011101110","0000101001011010010110100101","0000011100110111001101110011","0000010000110100001101000011","0000100100001001000010010000","0000110010111100101111001011","0000110010001100100011001000","0000110111111101111111011111","0000111111001111110011111100","0000100111011001110110011101","0000111011001110110011101100","0000110101101101011011010110","0000101101011011010110110101","0000011001010110010101100101","0000011011110110111101101111","0001000000000000000000000000","0000100111011001110110011101","0000101101101011011010110110","0000011110010111100101111001","0000101110011011100110111001","0000100110001001100010011000","0000100000101000001010000010","0000011000100110001001100010","0000001001010010010100100101","0000011010010110100101101001","0000001111100011111000111110","0000010001100100011001000110","0001000000000000000000000000","0001000000000000000000000000","0000010001000100010001000100","0000010011010100110101001101","0000001011110010111100101111","0000000011110000111100001111","0000010001000100010001000100","0000001101010011010100110101","0000001111100011111000111110","0000000001000000010000000100","0000010001010100010101000101","0000100111101001111010011110","0000111010011110100111101001","0000110010011100100111001001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111011111110111111101111","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000111111111111111111111111","0000111101001111010011110100","0000111100001111000011110000","0000111110001111100011111000","0000101011101010111010101110","0000000110100001101000011010","0000100011101000111010001110","0000111110011111100111111001","0000111111001111110011111100","0000111101011111010111110101","0000111110001111100011111000","0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000110111111101111111011111","0000110100111101001111010011","0000101110001011100010111000","0000110010011100100111001001","0000110110101101101011011010","0000110010011100100111001001","0000111110101111101011111010","0000111000101110001011100010","0000101100111011001110110011","0000110001011100010111000101","0000101110101011101010111010","0000011011100110111001101110","0000011111010111110101111101","0000101101101011011010110110","0000011111010111110101111101","0000011010100110101001101010","0000010101010101010101010101","0000100010011000100110001001","0000010110110101101101011011","0000110111001101110011011100","0000011100110111001101110011","0000010000000100000001000000","0000001111000011110000111100","0000100110001001100010011000","0000111010101110101011101010","0000110011011100110111001101","0000100010001000100010001000","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111011111110111111101","0000111111001111110011111100","0000111111001111110011111100","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111101011111010111110101","0000111111111111111111111111","0000110000101100001011000010","0000111100111111001111110011","0000110010001100100011001000","0000011110100111101001111010","0000111011111110111111101111","0000111101011111010111110101","0000111100111111001111110011","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111011111110111111101111","0000111111111111111111111111","0000111101111111011111110111","0000111010011110100111101001","0000110001011100010111000101","0000001111110011111100111111","0000000000100000001000000010","0000001100010011000100110001","0000111100011111000111110001","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111100001111000011110000","0000110011001100110011001100","0001000000000000000000000000","0000011100100111001001110010","0000100001101000011010000110","0000011010010110100101101001","0000101010101010101010101010","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000110000011100000111000001","0000101111101011111010111110","0000111001011110010111100101","0000100101011001010110010101","0000111000011110000111100001","0000111111111111111111111111","0000111011001110110011101100","0000111101101111011011110110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110000001100000011000000","0000110101001101010011010100","0000111111111111111111111111","0000111110011111100111111001","0000101011111010111110101111","0000100001001000010010000100","0000011001010110010101100101","0000010101010101010101010101","0000011110010111100101111001","0000010010100100101001001010","0000010111010101110101011101","0000101010011010100110101001","0000100100111001001110010011","0000111010101110101011101010","0000111110011111100111111001","0000111010011110100111101001","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111101101111011011110110","0000111110101111101011111010","0000111100111111001111110011","0000111101011111010111110101","0000111111111111111111111111","0000111111101111111011111110","0000111100101111001011110010","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000100010001000100010001000","0000010101110101011101010111","0001000000000000000000000000","0000011111000111110001111100","0000100101101001011010010110","0000100001111000011110000111","0000110110101101101011011010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111000111110001111100011","0000111000001110000011100000","0000100011011000110110001101","0000001010110010101100101011","0000010101100101011001010110","0000011100000111000001110000","0000100001001000010010000100","0000101000111010001110100011","0000110010001100100011001000","0000101101111011011110110111","0000111000101110001011100010","0000100100101001001010010010","0000101110001011100010111000","0000100001101000011010000110","0000101011111010111110101111","0000000011100000111000001110","0000010001000100010001000100","0000011111010111110101111101","0000011111010111110101111101","0000100110101001101010011010","0000110110111101101111011011","0000111111111111111111111111","0000101110101011101010111010","0000101111101011111010111110","0000011111000111110001111100","0000001100010011000100110001","0000000001010000010100000101","0000000110100001101000011010","0000000111100001111000011110","0000010010110100101101001011","0000011010000110100001101000","0000010000100100001001000010","0001000000000000000000000000","0000011011100110111001101110","0000101011111010111110101111","0000000100010001000100010001","0000001000010010000100100001","0000001011100010111000101110","0000001110010011100100111001","0000101000011010000110100001","0000100110111001101110011011","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110011111100111111001","0000111111001111110011111100","0000111110011111100111111001","0000111110101111101011111010","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000110110001101100011011000","0000010110100101101001011010","0000100100011001000110010001","0000111111111111111111111111","0000111010011110100111101001","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111000001110000011100000","0000110011111100111111001111","0000110001001100010011000100","0000111100111111001111110011","0000111011011110110111101101","0000111111111111111111111111","0000111001101110011011100110","0000111101111111011111110111","0000111111111111111111111111","0000111000001110000011100000","0000111001101110011011100110","0000101001001010010010100100","0000100000011000000110000001","0000100000011000000110000001","0000101110011011100110111001","0000010011010100110101001101","0000101010111010101110101011","0000011100110111001101110011","0000101100101011001010110010","0000010011000100110001001100","0000011100110111001101110011","0000010010100100101001001010","0000101010001010100010101000","0000110001001100010011000100","0000111111111111111111111111","0000010110110101101101011011","0000111110001111100011111000","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111110011111100111111001","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000101111001011110010111100","0000111010101110101011101010","0000101101001011010010110100","0000100101111001011110010111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111011111110111111101","0000111100011111000111110001","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111100101111001011110010","0000110000001100000011000000","0000010100110101001101010011","0001000000000000000000000000","0000011110110111101101111011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111101001111010011110100","0000111110001111100011111000","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000001000010010000100100001","0000011011010110110101101101","0000100000001000000010000000","0000100011111000111110001111","0000011100100111001001110010","0000110111101101111011011110","0000111110111111101111111011","0000111111111111111111111111","0000100101111001011110010111","0000100101001001010010010100","0000110010101100101011001010","0000101110001011100010111000","0000110110001101100011011000","0000111111111111111111111111","0000111101001111010011110100","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000110001001100010011000100","0000111110111111101111111011","0000111111111111111111111111","0000100101001001010010010100","0000101011011010110110101101","0000011101110111011101110111","0000010101010101010101010101","0000001000110010001100100011","0000100101101001011010010110","0000001010110010101100101011","0000100111011001110110011101","0000111101001111010011110100","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111011101110111011101110","0000111101001111010011110100","0000111110101111101011111010","0000111100001111000011110000","0000111111111111111111111111","0000111101111111011111110111","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111110101111101011111010","0000111010001110100011101000","0000100010111000101110001011","0000011101100111011001110110","0000000111000001110000011100","0000001111010011110100111101","0000110110111101101111011011","0000011011100110111001101110","0000101000111010001110100011","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111000101110001011100010","0000011010010110100101101001","0000001101110011011100110111","0000010010100100101001001010","0000010100100101001001010010","0000011101000111010001110100","0000101111011011110110111101","0000101101001011010010110100","0000100101011001010110010101","0000110111011101110111011101","0000011111110111111101111111","0000100001001000010010000100","0000011001110110011101100111","0000010101110101011101010111","0000000001000000010000000100","0000001011000010110000101100","0000010110110101101101011011","0000011001010110010101100101","0000011000110110001101100011","0000101010001010100010101000","0000101101011011010110110101","0000011101110111011101110111","0000001001100010011000100110","0000000011000000110000001100","0000010100010101000101010001","0000001111110011111100111111","0000010110100101101001011010","0000001110100011101000111010","0000010110010101100101011001","0000001100010011000100110001","0000000000100000001000000010","0000001011000010110000101100","0000011010100110101001101010","0000010000010100000101000001","0001000000000000000000000000","0000011001100110011001100110","0000011100000111000001110000","0000100010111000101110001011","0000101110001011100010111000","0000101101111011011110110111","0000111010001110100011101000","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000100011101000111010001110","0000011101100111011001110110","0000111001011110010111100101","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000111101101111011011110110","0000111011111110111111101111","0000111100011111000111110001","0000111111111111111111111111","0000111010111110101111101011","0000111000111110001111100011","0000110001111100011111000111","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111101111111011111110","0000111101101111011011110110","0000111110101111101011111010","0000111101011111010111110101","0000101010001010100010101000","0000100101011001010110010101","0000101001011010010110100101","0000010111110101111101011111","0000100000111000001110000011","0000011010010110100101101001","0000100100001001000010010000","0000010001000100010001000100","0000011111010111110101111101","0000101100001011000010110000","0000100000011000000110000001","0000100110111001101110011011","0000110101101101011011010110","0000101001111010011110100111","0000101111111011111110111111","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111110001111100011111000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111011111110111111101","0000111110011111100111111001","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000110001001100010011000100","0000111111111111111111111111","0000100101111001011110010111","0000110100101101001011010010","0000111111001111110011111100","0000111011111110111111101111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111100001111000011110000","0000110001111100011111000111","0000001010110010101100101011","0000000001000000010000000100","0000110000101100001011000010","0000111101001111010011110100","0000111111011111110111111101","0000111100111111001111110011","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111101111111011111110","0000111110011111100111111001","0000111101111111011111110111","0000111110011111100111111001","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000100101011001010110010101","0000001000100010001000100010","0000101000111010001110100011","0000011111100111111001111110","0000100110111001101110011011","0000100101101001011010010110","0000110111011101110111011101","0000111011011110110111101101","0000010111100101111001011110","0000011011010110110101101101","0000101010111010101110101011","0000110100101101001011010010","0000110100111101001111010011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000110100011101000111010001","0000111101111111011111110111","0000111110011111100111111001","0000100100111001001110010011","0000100000011000000110000001","0000011100110111001101110011","0000001111000011110000111100","0000010110000101100001011000","0000010100110101001101010011","0000100100101001001010010010","0000101011011010110110101101","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000011001100110011001100110","0000011011110110111101101111","0000011010110110101101101011","0001000000000000000000000000","0000111001011110010111100101","0000110000011100000111000001","0000011110100111101001111010","0000110100001101000011010000","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000101100101011001010110010","0000001011110010111100101111","0000011100100111001001110010","0000011100010111000101110001","0000010000110100001101000011","0000011011110110111101101111","0000100010101000101010001010","0000010010100100101001001010","0000101010011010100110101001","0000100100111001001110010011","0000011111000111110001111100","0000011101100111011001110110","0000100010111000101110001011","0000001011000010110000101100","0000000011110000111100001111","0000000000100000001000000010","0000010011000100110001001100","0000001011100010111000101110","0000010000110100001101000011","0000001010010010100100101001","0000001000110010001100100011","0000001110000011100000111000","0000011111010111110101111101","0000100010001000100010001000","0000001011010010110100101101","0000010001000100010001000100","0000000111010001110100011101","0000011110010111100101111001","0000000110110001101100011011","0000000010110000101100001011","0000011001000110010001100100","0000011111010111110101111101","0000011011110110111101101111","0000010101110101011101010111","0000001000100010001000100010","0000011111000111110001111100","0000010111000101110001011100","0000101001011010010110100101","0000101000111010001110100011","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111010111110101111101011","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000100011011000110110001101","0000110011101100111011001110","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111001001110010011100100","0000111011001110110011101100","0000110001001100010011000100","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111001101110011011100110","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000110101001101010011010100","0000101100001011000010110000","0000100101001001010010010100","0000100000111000001110000011","0000011001110110011101100111","0000011100100111001001110010","0000011010100110101001101010","0000001101100011011000110110","0000011111010111110101111101","0000110011011100110111001101","0000100110001001100010011000","0000101001011010010110100101","0000110011011100110111001101","0000100000011000000110000001","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110101111101011111010","0000111110111111101111111011","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111011111110111111101111","0000101000101010001010100010","0000111001011110010111100101","0000111101101111011011110110","0000111111111111111111111111","0000111011111110111111101111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111101111111011111110","0000111110001111100011111000","0000111011111110111111101111","0000110001101100011011000110","0001000000000000000000000000","0000000101010001010100010101","0000110101101101011011010110","0000111101101111011011110110","0000111100011111000111110001","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111011011110110111101101","0000111110101111101011111010","0000111110101111101011111010","0000110111101101111011011110","0001000000000000000000000000","0000011100100111001001110010","0000101101101011011010110110","0000101011011010110110101101","0000101111111011111110111111","0000100110001001100010011000","0000110110101101101011011010","0000001110100011101000111010","0000011100110111001101110011","0000011101000111010001110100","0000101011011010110110101101","0000111100101111001011110010","0000111111111111111111111111","0000111100011111000111110001","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111101011111010111110101","0000111101001111010011110100","0000111110001111100011111000","0000110010011100100111001001","0000101111001011110010111100","0000011111110111111101111111","0000011001010110010101100101","0001000000000000000000000000","0000010101100101011001010110","0000011000100110001001100010","0000011100110111001101110011","0000111111001111110011111100","0000111110011111100111111001","0000111100011111000111110001","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000101110111011101110111011","0000011001000110010001100100","0000010100010101000101010001","0000101100011011000110110001","0000000100110001001100010011","0000011010000110100001101000","0000111011101110111011101110","0000011111110111111101111111","0000101000011010000110100001","0000110110011101100111011001","0000111100101111001011110010","0000111100011111000111110001","0000111111101111111011111110","0000111010111110101111101011","0000111100101111001011110010","0000111111111111111111111111","0000111100011111000111110001","0000100101111001011110010111","0000001010100010101000101010","0000001011010010110100101101","0000011000010110000101100001","0000011001010110010101100101","0000011010110110101101101011","0000011011100110111001101110","0000100010111000101110001011","0000101000101010001010100010","0000011011110110111101101111","0000001111100011111000111110","0000010011110100111101001111","0000011101100111011001110110","0000001100100011001000110010","0000000101010001010100010101","0000000101110001011100010111","0001000000000000000000000000","0000000001100000011000000110","0001000000000000000000000000","0000001000000010000000100000","0000001010100010101000101010","0000010111010101110101011101","0000010100010101000101010001","0000001100110011001100110011","0000001100010011000100110001","0000001001010010010100100101","0000010100000101000001010000","0000000001100000011000000110","0000001110010011100100111001","0000011000010110000101100001","0000001100000011000000110000","0000011001110110011101100111","0000010101010101010101010101","0000011000010110000101100001","0000000010110000101100001011","0000001010010010100100101001","0000001111000011110000111100","0000101110011011100110111001","0000011101110111011101110111","0000111101101111011011110110","0000111100011111000111110001","0000111111101111111011111110","0000111110111111101111111011","0000111011001110110011101100","0000101010101010101010101010","0000111101111111011111110111","0000111110111111101111111011","0000111110011111100111111001","0000111011001110110011101100","0000111011101110111011101110","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111100111111001111110011","0000111010011110100111101001","0000110111001101110011011100","0000111011001110110011101100","0000111011111110111111101111","0000101111001011110010111100","0000111001011110010111100101","0000111011011110110111101101","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111011101110111011101110","0000101001011010010110100101","0000011110010111100101111001","0000010110000101100001011000","0000011001100110011001100110","0000011001010110010101100101","0000010010110100101101001011","0000011011010110110101101101","0000100100011001000110010001","0000110001011100010111000101","0000011010110110101101101011","0000100110111001101110011011","0000101111111011111110111111","0000100001101000011010000110","0000111101101111011011110110","0000111101111111011111110111","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111100101111001011110010","0000111111011111110111111101","0000111100101111001011110010","0000111001011110010111100101","0000111110101111101011111010","0000111111111111111111111111","0000110110011101100111011001","0000110011001100110011001100","0000111100111111001111110011","0000110101101101011011010110","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111101101111011011110110","0000111101001111010011110100","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000011111010111110101111101","0000000111100001111000011110","0000010000000100000001000000","0000111010011110100111101001","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111011111110111111101111","0000111111111111111111111111","0000111101101111011011110110","0000111011011110110111101101","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111011001110110011101100","0000001000100010001000100010","0000000010110000101100001011","0000100001001000010010000100","0000101100001011000010110000","0000110000111100001111000011","0000111010101110101011101010","0000011100100111001001110010","0000000000010000000100000001","0000011010100110101001101010","0000011001110110011101100111","0000100110001001100010011000","0000111101001111010011110100","0000111100111111001111110011","0000111101111111011111110111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111001111110011111100","0000111011101110111011101110","0000111011101110111011101110","0000111111111111111111111111","0000111111001111110011111100","0000100100101001001010010010","0000111011011110110111101101","0000100000001000000010000000","0000001110110011101100111011","0000000101000001010000010100","0000011110000111100001111000","0000010011010100110101001101","0000100110111001101110011011","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111100011111000111110001","0000111111111111111111111111","0000111111101111111011111110","0000110111101101111011011110","0000101010001010100010101000","0000010100110101001101010011","0000001001000010010000100100","0000011000000110000001100000","0000011100010111000101110001","0000100100011001000110010001","0001000000000000000000000000","0000010000100100001001000010","0000101000011010000110100001","0000001001100010011000100110","0000011110010111100101111001","0000110101001101010011010100","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000101110011011100110111001","0000101111101011111010111110","0000011111110111111101111111","0000001100110011001100110011","0000000101000001010000010100","0001000000000000000000000000","0000001001100010011000100110","0000010100000101000001010000","0000010010110100101101001011","0000011110100111101001111010","0000011110110111101101111011","0000010010100100101001001010","0000010000000100000001000000","0000001010000010100000101000","0000001111000011110000111100","0000010111110101111101011111","0000011101100111011001110110","0000001111100011111000111110","0000001101000011010000110100","0000001011010010110100101101","0001000000000000000000000000","0000001010010010100100101001","0000001110000011100000111000","0001000000000000000000000000","0000001001010010010100100101","0000001000000010000000100000","0000001000000010000000100000","0000000010100000101000001010","0000001010000010100000101000","0000001111110011111100111111","0000001101100011011000110110","0000010111100101111001011110","0000011001000110010001100100","0000100110111001101110011011","0000010000110100001101000011","0000000001000000010000000100","0001000000000000000000000000","0000001100000011000000110000","0000110010011100100111001001","0000101101001011010010110100","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111001011110010111100101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111101111111011111110","0000111111101111111011111110","0000111100111111001111110011","0000110011001100110011001100","0000101111001011110010111100","0000111010011110100111101001","0000111111111111111111111111","0000011111010111110101111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111111011111110111111101","0000111000101110001011100010","0000101111111011111110111111","0000011100100111001001110010","0000100000001000000010000000","0000010110010101100101011001","0000010011110100111101001111","0000100101101001011010010110","0000010010000100100001001000","0000011100110111001101110011","0000011111010111110101111101","0000101000001010000010100000","0000100101001001010010010100","0000110001101100011011000110","0000100100001001000010010000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111010111110101111101011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111110101111101011111010","0000101110011011100110111001","0000111101101111011011110110","0000111111111111111111111111","0000101010101010101010101010","0000111101001111010011110100","0000110111011101110111011101","0000111000011110000111100001","0000111111011111110111111101","0000111011101110111011101110","0000111001111110011111100111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000000110110001101100011011","0000011010100110101001101010","0000011011010110110101101101","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101001111010011110100","0000111011101110111011101110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000010000100100001001000010","0001000000000000000000000000","0000010100000101000001010000","0000100111111001111110011111","0000111111111111111111111111","0000110010111100101111001011","0000001010010010100100101001","0000011000000110000001100000","0000010100110101001101010011","0000000101110001011100010111","0000110001011100010111000101","0000111010111110101111101011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110111001101110011011100","0000101110111011101110111011","0000110000001100000011000000","0000011011010110110101101101","0000000011010000110100001101","0000001011000010110000101100","0000011101100111011001110110","0000010000110100001101000011","0000101011101010111010101110","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000110101001101010011010100","0000101001101010011010100110","0000101011001010110010101100","0000111000101110001011100010","0000100001011000010110000101","0000001100010011000100110001","0000011000000110000001100000","0000100010111000101110001011","0000011100100111001001110010","0000010001100100011001000110","0000010001010100010101000101","0000011000000110000001100000","0000100111001001110010011100","0000100001001000010010000100","0000101011101010111010101110","0000100110001001100010011000","0000110010011100100111001001","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000101110001011100010111000","0000110100001101000011010000","0000101010001010100010101000","0000100111001001110010011100","0001000000000000000000000000","0000000000110000001100000011","0001000000000000000000000000","0000001101110011011100110111","0000001010100010101000101010","0000001001110010011100100111","0000001101010011010100110101","0000010101110101011101010111","0000100000101000001010000010","0000010110100101101001011010","0000011010000110100001101000","0000011111010111110101111101","0000100101001001010010010100","0000011011100110111001101110","0000100000111000001110000011","0000011100100111001001110010","0000010001010100010101000101","0000001000010010000100100001","0000010110100101101001011010","0000010011010100110101001101","0000000111110001111100011111","0001000000000000000000000000","0000001000000010000000100000","0000010000000100000001000000","0000001011100010111000101110","0000010011110100111101001111","0000100000011000000110000001","0000101010011010100110101001","0000101010001010100010101000","0000001111010011110100111101","0000000000010000000100000001","0000001011110010111100101111","0000010110110101101101011011","0000110100101101001011010010","0000101011011010110110101101","0000111100001111000011110000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100101111001011110010","0000111011101110111011101110","0000101000011010000110100001","0000111110011111100111111001","0000111100101111001011110010","0000100111111001111110011111","0000111000011110000111100001","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111001011110010111100101","0000100111011001110110011101","0000011100010111000101110001","0000010011110100111101001111","0000001010100010101000101010","0000011100100111001001110010","0000100000001000000010000000","0000010111110101111101011111","0000010110100101101001011010","0000110001111100011111000111","0000101010001010100010101000","0000101001111010011110100111","0000100111111001111110011111","0000110001011100010111000101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111011011110110111101101","0000111110111111101111111011","0000111101011111010111110101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000110100011101000111010001","0000111100101111001011110010","0000110010001100100011001000","0000110111101101111011011110","0000111111111111111111111111","0000101010011010100110101001","0000111100001111000011110000","0000111111111111111111111111","0000110101111101011111010111","0000111111111111111111111111","0000111100101111001011110010","0000111011111110111111101111","0000111111111111111111111111","0000101100011011000110110001","0000001000100010001000100010","0000011011010110110101101101","0000110010011100100111001001","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000011100010111000101110001","0000000001110000011100000111","0000000100100001001000010010","0000000001110000011100000111","0000101010001010100010101000","0000000110010001100100011001","0000010111000101110001011100","0000101110111011101110111011","0000010010000100100001001000","0000010111110101111101011111","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110111111101111111011","0000111110101111101011111010","0000110011011100110111001101","0000111011111110111111101111","0000011111000111110001111100","0000001011100010111000101110","0001000000000000000000000000","0000001100110011001100110011","0000011010000110100001101000","0000010001100100011001000110","0000101111111011111110111111","0000111010101110101011101010","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111011111110111111101111","0000110111011101110111011101","0000111001011110010111100101","0000111100111111001111110011","0000111111001111110011111100","0000110111111101111111011111","0000010111100101111001011110","0000010010000100100001001000","0000010001100100011001000110","0000100100101001001010010010","0000100000101000001010000010","0000011110010111100101111001","0000010001000100010001000100","0000010111100101111001011110","0000100100111001001110010011","0000100101001001010010010100","0000011100010111000101110001","0000110010011100100111001001","0000101001111010011110100111","0000011010100110101001101010","0000100111101001111010011110","0000111010101110101011101010","0000111101011111010111110101","0000111101011111010111110101","0000111000101110001011100010","0000111000111110001111100011","0000110000111100001111000011","0000111010001110100011101000","0000111110101111101011111010","0000011111010111110101111101","0000010100100101001001010010","0000010110000101100001011000","0000010100010101000101010001","0000010101110101011101010111","0000011110000111100001111000","0000100110101001101010011010","0000101010111010101110101011","0000101110011011100110111001","0000110000001100000011000000","0000111011001110110011101100","0000111010011110100111101001","0000111011001110110011101100","0000110101001101010011010100","0000001111000011110000111100","0000100000101000001010000010","0000010010000100100001001000","0000010001000100010001000100","0000011011000110110001101100","0000100000011000000110000001","0000010010000100100001001000","0000000111100001111000011110","0000000010010000100100001001","0000001001010010010100100101","0000001001000010010000100100","0000001011100010111000101110","0000011100110111001101110011","0000100111011001110110011101","0000101011001010110010101100","0000010111100101111001011110","0000000010010000100100001001","0001000000000000000000000000","0000100010101000101010001010","0000010000100100001001000010","0000101100011011000110110001","0000100111011001110110011101","0000110010101100101011001010","0000111101111111011111110111","0000111011001110110011101100","0000111111111111111111111111","0000111001001110010011100100","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101101111011011110110","0000101010111010101110101011","0000111110101111101011111010","0000111101011111010111110101","0000111010011110100111101001","0000101011101010111010101110","0000111010111110101111101011","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000110100101101001011010010","0000100101111001011110010111","0000011101110111011101110111","0000010111010101110101011101","0000011101000111010001110100","0000011011010110110101101101","0000011010000110100001101000","0000010101010101010101010101","0000100011111000111110001111","0000101111001011110010111100","0000100111101001111010011110","0000100110101001101010011010","0000101010101010101010101010","0000110010101100101011001010","0000111100111111001111110011","0000111110111111101111111011","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111110011111100111111001","0000111110111111101111111011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000110100101101001011010010","0000111111111111111111111111","0000111011011110110111101101","0000111001101110011011100110","0000111101001111010011110100","0000110100111101001111010011","0000111010111110101111101011","0000111100111111001111110011","0000111000001110000011100000","0000110110001101100011011000","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0001000000000000000000000000","0000011101110111011101110111","0000001101100011011000110110","0000110101101101011011010110","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000100011011000110110001101","0000000100100001001000010010","0000000011010000110100001101","0000001011110010111100101111","0000000111110001111100011111","0000010010010100100101001001","0000101110011011100110111001","0000011100100111001001110010","0000011100010111000101110001","0000110000111100001111000011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111011111110111111101111","0000110010101100101011001010","0000110011011100110111001101","0000100001011000010110000101","0000000100000001000000010000","0000001101100011011000110110","0000011011000110110001101100","0000010100110101001101010011","0000011110100111101001111010","0000110000111100001111000011","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111011111110111111101","0000111101001111010011110100","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000101111001011110010111100","0000010111110101111101011111","0000011110010111100101111001","0000011000100110001001100010","0000100010101000101010001010","0000001100100011001000110010","0000001110110011101100111011","0000000110110001101100011011","0000000110000001100000011000","0000000011110000111100001111","0000010101010101010101010101","0000101001011010010110100101","0000111000111110001111100011","0000110010101100101011001010","0000011111110111111101111111","0000101101101011011010110110","0000111001011110010111100101","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111100101111001011110010","0000110111011101110111011101","0000110010101100101011001010","0000101010101010101010101010","0000110110011101100111011001","0000011110100111101001111010","0000001110100011101000111010","0000011010010110100101101001","0000101000011010000110100001","0000100011101000111010001110","0000101010001010100010101000","0000111101101111011011110110","0000111111101111111011111110","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000100111111001111110011111","0000010111100101111001011110","0000010101110101011101010111","0000001111110011111100111111","0000010101100101011001010110","0000100100111001001110010011","0000000110110001101100011011","0000000010010000100100001001","0001000000000000000000000000","0000001110000011100000111000","0000001011010010110100101101","0000011000110110001101100011","0000110010101100101011001010","0000110001111100011111000111","0000100101101001011010010110","0000110000101100001011000010","0000010111100101111001011110","0000000010110000101100001011","0000000011110000111100001111","0000100001001000010010000100","0000010000110100001101000011","0000011111000111110001111100","0000110001011100010111000101","0000110001101100011011000110","0000111111111111111111111111","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000101110111011101110111011","0000100110101001101010011010","0000010001100100011001000110","0000100111101001111010011110","0000110111011101110111011101","0000111001001110010011100100","0000110010101100101011001010","0000111100111111001111110011","0000110111101101111011011110","0000111110001111100011111000","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111101011111010111110101","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000101101101011011010110110","0000100100001001000010010000","0000011011010110110101101101","0000101001101010011010100110","0000010101100101011001010110","0000100001101000011010000110","0000010100000101000001010000","0000100001011000010110000101","0000100110011001100110011001","0000110100001101000011010000","0000100001111000011110000111","0000101001001010010010100100","0000110011111100111111001111","0000101110001011100010111000","0000101111111011111110111111","0000111011101110111011101110","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000111100101111001011110010","0000111011011110110111101101","0000111101101111011011110110","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000110111101101111011011110","0000110100001101000011010000","0000111011111110111111101111","0000111011101110111011101110","0000110110111101101111011011","0000111000111110001111100011","0000111011111110111111101111","0000110111011101110111011101","0000111010001110100011101000","0000111101011111010111110101","0000110100101101001011010010","0000111111111111111111111111","0000111100111111001111110011","0000011111100111111001111110","0000001100010011000100110001","0000101010011010100110101001","0000001000100010001000100010","0000111010011110100111101001","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110000011100000111000001","0000000010000000100000001000","0000001000000010000000100000","0000010101100101011001010110","0000011011000110110001101100","0000011011010110110101101101","0000001101010011010100110101","0000010001000100010001000100","0000010111000101110001011100","0000101011011010110110101101","0000110011011100110111001101","0000111010101110101011101010","0000111011111110111111101111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000111010101110101011101010","0000100000001000000010000000","0000110001011100010111000101","0001000000000000000000000000","0000100010001000100010001000","0000011101000111010001110100","0000010110100101101001011010","0000011101000111010001110100","0000101111001011110010111100","0000111111001111110011111100","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101001111010011110100","0000111101101111011011110110","0000101101111011011110110111","0000100010001000100010001000","0000100010001000100010001000","0000101100101011001010110010","0000110100111101001111010011","0000011111000111110001111100","0000110000011100000111000001","0000111011011110110111101101","0000101110001011100010111000","0000011101010111010101110101","0000001100010011000100110001","0000010101000101010001010100","0000100010111000101110001011","0000110111111101111111011111","0000111101101111011011110110","0000011111100111111001111110","0000101001011010010110100101","0000111010101110101011101010","0000111100111111001111110011","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000110101111101011111010111","0000110011111100111111001111","0000100111101001111010011110","0000100000101000001010000010","0000101011111010111110101111","0000110100111101001111010011","0000110111111101111111011111","0000110011011100110111001101","0000101001101010011010100110","0000110000001100000011000000","0000110000111100001111000011","0000110101111101011111010111","0000111100101111001011110010","0000111000011110000111100001","0000110110101101101011011010","0000011001010110010101100101","0000011000010110000101100001","0000010001100100011001000110","0000010101100101011001010110","0000011001010110010101100101","0000001000000010000000100000","0000000010010000100100001001","0000000111110001111100011111","0000010001000100010001000100","0000011010100110101001101010","0000101000111010001110100011","0000110010001100100011001000","0000100001011000010110000101","0000100111111001111110011111","0000101010101010101010101010","0000101000001010000010100000","0000011100100111001001110010","0000000110100001101000011010","0000000010010000100100001001","0000011100100111001001110010","0000100011011000110110001101","0000010110100101101001011010","0000010011110100111101001111","0000011111010111110101111101","0000101010101010101010101010","0000110011001100110011001100","0000101101011011010110110101","0000100011011000110110001101","0000010011000100110001001100","0000010110010101100101011001","0000010001010100010101000101","0000001101010011010100110101","0000110000111100001111000011","0000110010101100101011001010","0000101001111010011110100111","0000110111001101110011011100","0000111000001110000011100000","0000111110111111101111111011","0000111111101111111011111110","0000111011001110110011101100","0000111111001111110011111100","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000101010001010100010101000","0000100011001000110010001100","0000011111110111111101111111","0000101001011010010110100101","0000001110110011101100111011","0000011110100111101001111010","0000100101001001010010010100","0000011110010111100101111001","0000100101111001011110010111","0000101010011010100110101001","0000101001011010010110100101","0000101000101010001010100010","0000101111101011111010111110","0000100010001000100010001000","0000011101000111010001110100","0000100010111000101110001011","0000110111011101110111011101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111110011111100111111001","0000111100101111001011110010","0000111100101111001011110010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000110100011101000111010001","0000110100001101000011010000","0000110001111100011111000111","0000110100111101001111010011","0000110010011100100111001001","0000110110001101100011011000","0000110101101101011011010110","0000110000111100001111000011","0000111000101110001011100010","0000101110001011100010111000","0000110101101101011011010110","0000111011001110110011101100","0000101110111011101110111011","0000000000110000001100000011","0000101011111010111110101111","0000000101000001010000010100","0000100000101000001010000010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0001000000000000000000000000","0000011110110111101101111011","0000010010010100100101001001","0000010110000101100001011000","0000011101100111011001110110","0000010110110101101101011011","0000010111010101110101011101","0000110011011100110111001101","0000111000101110001011100010","0000111011101110111011101110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111101001111010011110100","0000111100011111000111110001","0000111000101110001011100010","0000100101011001010110010101","0000110011101100111011001110","0000000010010000100100001001","0000100101111001011110010111","0000101011011010110110101101","0000010110100101101001011010","0000100011001000110010001100","0000100011101000111010001110","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000110011111100111111001111","0000110101011101010111010101","0000110011111100111111001111","0000111100001111000011110000","0000110101111101011111010111","0000011011000110110001101100","0000110100111101001111010011","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111110111111101111111011","0000101110111011101110111011","0000100100001001000010010000","0000011101010111010101110101","0000011001100110011001100110","0000110101111101011111010111","0000110001111100011111000111","0000011110010111100101111001","0000111111111111111111111111","0000111100101111001011110010","0000111101001111010011110100","0000111111111111111111111111","0000111011111110111111101111","0000111111011111110111111101","0000111101111111011111110111","0000111110111111101111111011","0000110111011101110111011101","0000110111001101110011011100","0000110111001101110011011100","0000110101011101010111010101","0000110110101101101011011010","0000111001001110010011100100","0000110111111101111111011111","0000110110011101100111011001","0000110101101101011011010110","0000111010011110100111101001","0000111001011110010111100101","0000111010111110101111101011","0000011101000111010001110100","0000110000001100000011000000","0000010110110101101101011011","0000100000001000000010000000","0000011010100110101001101010","0000001001000010010000100100","0000011100110111001101110011","0000001010100010101000101010","0000001000000010000000100000","0000000110010001100100011001","0000100101001001010010010100","0000011111000111110001111100","0000011111110111111101111111","0000011100000111000001110000","0000100111101001111010011110","0000101001101010011010100110","0000101111111011111110111111","0000100111111001111110011111","0000101000101010001010100010","0000000101000001010000010100","0001000000000000000000000000","0000001111010011110100111101","0000101011101010111010101110","0000101001101010011010100110","0000001110000011100000111000","0000010101100101011001010110","0000010101110101011101010111","0000010001110100011101000111","0000011000010110000101100001","0000011101110111011101110111","0000010101000101010001010100","0000010010000100100001001000","0000100101011001010110010101","0000100010111000101110001011","0000101001001010010010100100","0000111011011110110111101101","0000110101111101011111010111","0000111111111111111111111111","0000111010011110100111101001","0000111101101111011011110110","0000111111111111111111111111","0000111011011110110111101101","0000111110001111100011111000","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111001001110010011100100","0000101100111011001110110011","0000100100001001000010010000","0000100101001001010010010100","0000010100010101000101010001","0000011011000110110001101100","0000100000111000001110000011","0000100010011000100110001001","0000001110000011100000111000","0000100011111000111110001111","0000011100110111001101110011","0000100010101000101010001010","0000011101010111010101110101","0000100101001001010010010100","0000011100000111000001110000","0000010111100101111001011110","0000010011000100110001001100","0000110001001100010011000100","0000111010011110100111101001","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111101101111011011110110","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111010011110100111101001","0000110111101101111011011110","0000110001101100011011000110","0000101000101010001010100010","0000100110001001100010011000","0000101110111011101110111011","0000101101011011010110110101","0000110000111100001111000011","0000100111011001110110011101","0000101010011010100110101001","0000110100001101000011010000","0000101000011010000110100001","0000101010101010101010101010","0000110110001101100011011000","0000000000100000001000000010","0000100000011000000110000001","0000010110010101100101011001","0000000011100000111000001110","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000000101100001011000010110","0000011111110111111101111111","0000100000111000001110000011","0000100001111000011110000111","0000100011111000111110001111","0000100010011000100110001001","0000101100101011001010110010","0000100010001000100010001000","0000100011101000111010001110","0000110000001100000011000000","0000111011001110110011101100","0000111000011110000111100001","0000111110001111100011111000","0000111001101110011011100110","0000111100101111001011110010","0000111111011111110111111101","0000111100111111001111110011","0000111110011111100111111001","0000111111101111111011111110","0000111101001111010011110100","0000100001011000010110000101","0000111010101110101011101010","0000101000001010000010100000","0000010010110100101101001011","0000101000101010001010100010","0000110111011101110111011101","0000101010001010100010101000","0000100000011000000110000001","0000100011011000110110001101","0000101001111010011110100111","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111110111111101111111011","0000111111001111110011111100","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111100111111001111110011","0000111111111111111111111111","0000111101001111010011110100","0000110001101100011011000110","0000110010011100100111001001","0000111101011111010111110101","0000110110011101100111011001","0000111111011111110111111101","0000111010101110101011101010","0000100001101000011010000110","0000111011001110110011101100","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000110110001101100011011000","0000011101010111010101110101","0000000000010000000100000001","0000011010100110101001101010","0000110011011100110111001101","0000011011100110111001101110","0000110111101101111011011110","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000111011001110110011101100","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000110111101101111011011110","0000110100111101001111010011","0000110001011100010111000101","0000110000011100000111000001","0000111000111110001111100011","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000101111011011110110111101","0000110000111100001111000011","0000101010011010100110101001","0000011111010111110101111101","0000100101001001010010010100","0000011010110110101101101011","0000001100100011001000110010","0000011100100111001001110010","0000001011000010110000101100","0000000010110000101100001011","0000001100010011000100110001","0000100100101001001010010010","0000011100110111001101110011","0000001110100011101000111010","0000100001101000011010000110","0000011011000110110001101100","0000110011101100111011001110","0000111001101110011011100110","0000110101001101010011010100","0000101101011011010110110101","0000100110011001100110011001","0000101001001010010010100100","0000000110000001100000011000","0000000000100000001000000010","0000010001110100011101000111","0000011100000111000001110000","0000011000100110001001100010","0000010101110101011101010111","0000010010110100101101001011","0000001111100011111000111110","0000001001000010010000100100","0000000011010000110100001101","0000011111110111111101111111","0000100101111001011110010111","0000101111101011111010111110","0000110001101100011011000110","0000101100111011001110110011","0000111111101111111011111110","0000111000011110000111100001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000110010111100101111001011","0000110010011100100111001001","0000101000011010000110100001","0000101010011010100110101001","0000010001100100011001000110","0000010101110101011101010111","0000010100100101001001010010","0000010111110101111101011111","0000011100100111001001110010","0000010111110101111101011111","0000011100110111001101110011","0000100000101000001010000010","0000010100010101000101010001","0000011100100111001001110010","0000011101010111010101110101","0000010101000101010001010100","0000000111110001111100011111","0000100110101001101010011010","0000110010011100100111001001","0000111001011110010111100101","0000111010001110100011101000","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100001111000011110000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110001011100010111000101","0000101101001011010010110100","0000101110101011101010111010","0000101101101011011010110110","0000011000000110000001100000","0000011011110110111101101111","0000101001101010011010100110","0000100110011001100110011001","0000101000101010001010100010","0000011111010111110101111101","0000100111111001111110011111","0000101110111011101110111011","0000100100011001000110010001","0000011011100110111001101110","0000000111010001110100011101","0000011000010110000101100001","0000101110001011100010111000","0000001011110010111100101111","0000011111000111110001111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000010100010101000101010001","0000010011010100110101001101","0000101011101010111010101110","0000101100111011001110110011","0000101101101011011010110110","0000101011011010110110101101","0000101101111011011110110111","0000111011011110110111101101","0000110101011101010111010101","0000110100001101000011010000","0000110011011100110111001101","0000101111101011111010111110","0000110100101101001011010010","0000110111011101110111011101","0000111101111111011111110111","0000111111101111111011111110","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000110001001100010011000100","0000011000110110001101100011","0000111111111111111111111111","0000010101010101010101010101","0000100001111000011110000111","0000100100111001001110010011","0000111111111111111111111111","0000110010101100101011001010","0000101000001010000010100000","0000100001111000011110000111","0000011101010111010101110101","0000101100011011000110110001","0000111100101111001011110010","0000111100111111001111110011","0000111101011111010111110101","0000111110001111100011111000","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111011111110111111101111","0000111111111111111111111111","0000111100111111001111110011","0000101111101011111010111110","0000110011001100110011001100","0000110011111100111111001111","0000111010011110100111101001","0000111111101111111011111110","0000111011011110110111101101","0000101111011011110110111101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111010001110100011101000","0000111101111111011111110111","0000110101011101010111010101","0000000100100001001000010010","0000000000010000000100000001","0000011101000111010001110100","0000100010111000101110001011","0000111000101110001011100010","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111011111110111111101111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111000111110001111100011","0000111000101110001011100010","0000110111001101110011011100","0000100101001001010010010100","0000011100100111001001110010","0000100111101001111010011110","0000010111110101111101011111","0000011000110110001101100011","0000001111100011111000111110","0000001000100010001000100010","0000000011100000111000001110","0000010110000101100001011000","0000011111110111111101111111","0000100110011001100110011001","0000000100010001000100010001","0000101101001011010010110100","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111100101111001011110010","0000110111111101111111011111","0000110000111100001111000011","0000101101001011010010110100","0000110111111101111111011111","0000011100110111001101110011","0000001110110011101100111011","0000000010010000100100001001","0000000001100000011000000110","0001000000000000000000000000","0001000000000000000000000000","0000000010010000100100001001","0000010000110100001101000011","0000100110011001100110011001","0000101100001011000010110000","0000100000001000000010000000","0000100111011001110110011101","0000110100001101000011010000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100011111000111110001","0000111011001110110011101100","0000110011101100111011001110","0000110100001101000011010000","0000101111011011110110111101","0000101001011010010110100101","0000010001100100011001000110","0000101010011010100110101001","0000100110101001101010011010","0000001001000010010000100100","0000011001110110011101100111","0000011111010111110101111101","0000011101000111010001110100","0000100110011001100110011001","0000110000101100001011000010","0000110110011101100111011001","0000011010110110101101101011","0000000000100000001000000010","0000010000100100001001000010","0000110000101100001011000010","0000110000011100000111000001","0000101000011010000110100001","0000101011001010110010101100","0000110101011101010111010101","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111100011111000111110001","0000111100111111001111110011","0000111100011111000111110001","0000110100111101001111010011","0000101011011010110110101101","0000101011011010110110101101","0000110001001100010011000100","0000110010111100101111001011","0000100100101001001010010010","0000100001111000011110000111","0000101000101010001010100010","0000100010001000100010001000","0000100010101000101010001010","0000100001011000010110000101","0000100011101000111010001110","0000100110111001101110011011","0000010011000100110001001100","0000000011010000110100001101","0000010000000100000001000000","0000110000001100000011000000","0000101011101010111010101110","0000000011010000110100001101","0000111000011110000111100001","0000111111101111111011111110","0000111110011111100111111001","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000011101000111010001110100","0001000000000000000000000000","0000110010011100100111001001","0000011111110111111101111111","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000110010111100101111001011","0000110100011101000111010001","0000110101001101010011010100","0000111001011110010111100101","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111100111111001111110011","0000011111110111111101111111","0000101001101010011010100110","0000111011111110111111101111","0000000010110000101100001011","0000101001001010010010100100","0000101001111010011110100111","0000111111111111111111111111","0000111111001111110011111100","0000110001101100011011000110","0000110000011100000111000001","0000100001111000011110000111","0000011101100111011001110110","0000111011001110110011101100","0000111011101110111011101110","0000111100011111000111110001","0000111101011111010111110101","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111011001110110011101100","0000110011001100110011001100","0000111011111110111111101111","0000110010101100101011001010","0000111111111111111111111111","0000111011111110111111101111","0000110000011100000111000001","0000110111011101110111011101","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000110111101101111011011110","0000110111001101110011011100","0000111010111110101111101011","0000011010010110100101101001","0000000000100000001000000010","0000000101000001010000010100","0000010010110100101101001011","0000111011101110111011101110","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111011011110110111101101","0000100010111000101110001011","0000011101100111011001110110","0000011110000111100001111000","0000101101001011010010110100","0000010000010100000101000001","0000010011010100110101001101","0000001010110010101100101011","0000000101010001010100010101","0000000001000000010000000100","0000000101010001010100010101","0000010100010101000101010001","0000011100010111000101110001","0000101010011010100110101001","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000110110111101101111011011","0000111100011111000111110001","0000111110001111100011111000","0000110111011101110111011101","0000111011011110110111101101","0000111111011111110111111101","0000101110101011101010111010","0000101111111011111110111111","0000101001011010010110100101","0000100100001001000010010000","0000100011101000111010001110","0000100101001001010010010100","0000101001011010010110100101","0000100101001001010010010100","0000101011101010111010101110","0000111001101110011011100110","0000111111111111111111111111","0000111011101110111011101110","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111110011111100111111001","0000111110111111101111111011","0000111111111111111111111111","0000110010111100101111001011","0000111000001110000011100000","0000110010101100101011001010","0000110101001101010011010100","0000100110011001100110011001","0000101101001011010010110100","0000101011111010111110101111","0000110000101100001011000010","0000100001011000010110000101","0000101000111010001110100011","0000001111100011111000111110","0000001111110011111100111111","0000011101100111011001110110","0000011101110111011101110111","0000101101111011011110110111","0000100111101001111010011110","0001000000000000000000000000","0000000000110000001100000011","0000011110010111100101111001","0000111100001111000011110000","0000111100001111000011110000","0000110000111100001111000011","0000100111011001110110011101","0000011111010111110101111101","0000011001110110011101100111","0000100000101000001010000010","0000101011101010111010101110","0000101111011011110110111101","0000110111001101110011011100","0000110011001100110011001100","0000110000001100000011000000","0000101100111011001110110011","0000101100111011001110110011","0000110101101101011011010110","0000111110111111101111111011","0000111111111111111111111111","0000101001011010010110100101","0000010111100101111001011110","0000010000100100001001000010","0000000110110001101100011011","0000000101000001010000010100","0000001001000010010000100100","0000000000010000000100000001","0000000001000000010000000100","0000000101100001011000010110","0000100000101000001010000010","0000110101001101010011010100","0000101100011011000110110001","0001000000000000000000000000","0000101011101010111010101110","0000111111001111110011111100","0000111111111111111111111111","0000111100111111001111110011","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000101010111010101110101011","0001000000000000000000000000","0000101111101011111010111110","0000101011101010111010101110","0000111111111111111111111111","0000111101101111011011110110","0000111100001111000011110000","0000110111101101111011011110","0000111100101111001011110010","0000111111111111111111111111","0000111110011111100111111001","0000111100011111000111110001","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111101101111011011110110","0000111111011111110111111101","0000110101001101010011010100","0000100001111000011110000111","0000110100011101000111010001","0000100110111001101110011011","0000000000010000000100000001","0000101000111010001110100011","0000110100111101001111010011","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000110011111100111111001111","0000111011111110111111101111","0000101010111010101110101011","0000011101110111011101110111","0000110110101101101011011010","0000111001101110011011100110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000110100101101001011010010","0000111111111111111111111111","0000111010001110100011101000","0000111100011111000111110001","0000111101111111011111110111","0000111001111110011111100111","0000110000101100001011000010","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111100111111001111110011","0000111100011111000111110001","0000110011001100110011001100","0000101100111011001110110011","0000110110011101100111011001","0000101001011010010110100101","0000010011100100111001001110","0001000000000000000000000000","0000000011000000110000001100","0000100100111001001110010011","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000110000101100001011000010","0000100010111000101110001011","0000011100110111001101110011","0000010101100101011001010110","0000000110000001100000011000","0000001110100011101000111010","0000010111010101110101011101","0000010011100100111001001110","0000000101110001011100010111","0000000011010000110100001101","0000010111110101111101011111","0000011100010111000101110001","0000011010100110101001101010","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000111010001110100011101000","0000101111111011111110111111","0000111111111111111111111111","0000111110011111100111111001","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111001111110011111100111","0000111011101110111011101110","0000111110101111101011111010","0000111111101111111011111110","0000111110101111101011111010","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111110111111101111111011","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111101101111011011110110","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000110100111101001111010011","0000110111001101110011011100","0000111100111111001111110011","0000111110101111101011111010","0000101000001010000010100000","0000110001001100010011000100","0000110100111101001111010011","0000101101011011010110110101","0000110010101100101011001010","0000101100001011000010110000","0000110011011100110111001101","0000110011111100111111001111","0000100100001001000010010000","0001000000000000000000000000","0000001000010010000100100001","0000100000101000001010000010","0000101001001010010010100100","0001000000000000000000000000","0000000100000001000000010000","0000101000011010000110100001","0000101010101010101010101010","0000101100111011001110110011","0000110100011101000111010001","0000111101001111010011110100","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000111111111111111111111111","0000110001101100011011000110","0000101111111011111110111111","0000101010001010100010101000","0000100101001001010010010100","0000101011111010111110101111","0000110010001100100011001000","0000011100000111000001110000","0000001010000010100000101000","0000001110100011101000111010","0000010100000101000001010000","0000011010110110101101101011","0000010111100101111001011110","0000010010100100101001001010","0000010000000100000001000000","0000000111100001111000011110","0000001101000011010000110100","0000010101010101010101010101","0000100101111001011110010111","0000110000001100000011000000","0000011100110111001101110011","0000001101110011011100110111","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000110001111100011111000111","0000000000010000000100000001","0000011010010110100101101001","0000101101011011010110110101","0000110110111101101111011011","0000111101111111011111110111","0000110111101101111011011110","0000100110001001100010011000","0000111111111111111111111111","0000111010011110100111101001","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111101001111010011110100","0000111110101111101011111010","0000111100101111001011110010","0000111110001111100011111000","0000110001001100010011000100","0000100011101000111010001110","0000101110101011101010111010","0000100011001000110010001100","0000000110110001101100011011","0000101101111011011110110111","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000111110001111100011","0000111110011111100111111001","0000110100011101000111010001","0000101011111010111110101111","0000110111011101110111011101","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111110101111101011111010","0000111111011111110111111101","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111100001111000011110000","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111001001110010011100100","0000110110011101100111011001","0000111110011111100111111001","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111110101111101011111010","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111110001111100011111000","0000111111001111110011111100","0000110111011101110111011101","0000101100001011000010110000","0000100101011001010110010101","0000100110001001100010011000","0000101111001011110010111100","0000100011111000111110001111","0000011101010111010101110101","0000001110110011101100111011","0000001001110010011100100111","0000101001101010011010100110","0000111100011111000111110001","0000111110011111100111111001","0000110111101101111011011110","0000111000101110001011100010","0000111110011111100111111001","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000110111101101111011011110","0000101011101010111010101110","0000010100110101001101010011","0000011101000111010001110100","0000011000000110000001100000","0000100001111000011110000111","0000001100010011000100110001","0000010110000101100001011000","0000011111100111111001111110","0000010101010101010101010101","0000001100000011000000110000","0000000100000001000000010000","0000001110110011101100111011","0000101100101011001010110010","0000100100001001000010010000","0000111111111111111111111111","0000111110001111100011111000","0000110001111100011111000111","0000111100001111000011110000","0000100100001001000010010000","0000111010101110101011101010","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111100111111001111110011","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000111010011110100111101001","0000111101111111011111110111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000110010101100101011001010","0000110100101101001011010010","0000111111111111111111111111","0000111011111110111111101111","0000110011101100111011001110","0000110001101100011011000110","0000110111101101111011011110","0000110001101100011011000110","0000110000011100000111000001","0000111001001110010011100100","0000111001001110010011100100","0000100101101001011010010110","0000111101001111010011110100","0000110100011101000111010001","0000101110001011100010111000","0000001000000010000000100000","0000001000100010001000100010","0000100000001000000010000000","0000001011000010110000101100","0001000000000000000000000000","0000100011111000111110001111","0000111001101110011011100110","0000101010011010100110101001","0000111110101111101011111010","0000110100011101000111010001","0000111000111110001111100011","0000111001001110010011100100","0000111001011110010111100101","0000111111111111111111111111","0000110110111101101111011011","0000011111100111111001111110","0000100101001001010010010100","0000010010010100100101001001","0000001010010010100100101001","0000000100010001000100010001","0000010111010101110101011101","0000100010011000100110001001","0000111010001110100011101000","0000110011101100111011001110","0000101100011011000110110001","0000100011101000111010001110","0000100010101000101010001010","0000001110100011101000111010","0000011011000110110001101100","0000011000100110001001100010","0000101011011010110110101101","0000100000101000001010000010","0000100101111001011110010111","0000100111011001110110011101","0000000001000000010000000100","0000111100011111000111110001","0000111111111111111111111111","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000001101000011010000110100","0000000001100000011000000110","0000101111101011111010111110","0000101001011010010110100101","0000111110111111101111111011","0000111000011110000111100001","0000101010101010101010101010","0000110000101100001011000010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000110000011100000111000001","0000100101101001011010010110","0000101010111010101110101011","0000100010011000100110001001","0000010010110100101101001011","0000100111001001110010011100","0000111111111111111111111111","0000111100111111001111110011","0000111100111111001111110011","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000111011001110110011101100","0000111111111111111111111111","0000100101111001011110010111","0000111101001111010011110100","0000111110011111100111111001","0000111101001111010011110100","0000111010011110100111101001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111011101110111011101110","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111101001111010011110100","0000111011111110111111101111","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111111101111111011111110","0000111101011111010111110101","0000111001011110010111100101","0000101101001011010010110100","0000011110100111101001111010","0000011100010111000101110001","0000100110111001101110011011","0000100010001000100010001000","0000100010001000100010001000","0000011001100110011001100110","0000000010000000100000001000","0000001101100011011000110110","0000011101110111011101110111","0000100110001001100010011000","0000100110111001101110011011","0000100100011001000110010001","0000100110011001100110011001","0000100110111001101110011011","0000101001111010011110100111","0000110010011100100111001001","0000101001011010010110100101","0000101011001010110010101100","0000010111000101110001011100","0000011010000110100001101000","0000001011000010110000101100","0000010100010101000101010001","0000010101000101010001010100","0000011111100111111001111110","0000100101001001010010010100","0000001101000011010000110100","0000101110011011100110111001","0000010100110101001101010011","0000000010010000100100001001","0000010011000100110001001100","0000100011101000111010001110","0000011101110111011101110111","0000110100111101001111010011","0000110010101100101011001010","0000110111011101110111011101","0000111010011110100111101001","0000101001001010010010100100","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111101001111010011110100","0000111010011110100111101001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111010001110100011101000","0000111111101111111011111110","0000111100011111000111110001","0000111001001110010011100100","0000111111111111111111111111","0000111100001111000011110000","0000110101011101010111010101","0000010101110101011101010111","0000111111111111111111111111","0000111001101110011011100110","0000110011111100111111001111","0000110001011100010111000101","0000111111111111111111111111","0000111000111110001111100011","0000101010111010101110101011","0000111110011111100111111001","0000111101111111011111110111","0000110110101101101011011010","0000110100001101000011010000","0000000001000000010000000100","0000000010100000101000001010","0000010010000100100001001000","0001000000000000000000000000","0000100001111000011110000111","0000110010001100100011001000","0000101000111010001110100011","0000101111011011110110111101","0000111111111111111111111111","0000111111101111111011111110","0000111011011110110111101101","0000111111111111111111111111","0000111111011111110111111101","0000100011001000110010001100","0000011011100110111001101110","0000001010100010101000101010","0000000110000001100000011000","0000010101100101011001010110","0000110000001100000011000000","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111000001110000011100000","0000101110001011100010111000","0000101001011010010110100101","0000101100011011000110110001","0000100010011000100110001001","0000101110001011100010111000","0000011111000111110001111100","0000011101100111011001110110","0000001100100011001000110010","0000100101011001010110010101","0000001001000010010000100100","0000101011101010111010101110","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000010111000101110001011100","0001000000000000000000000000","0000011000010110000101100001","0000101010011010100110101001","0000110010001100100011001000","0000111011001110110011101100","0000110001011100010111000101","0000110010111100101111001011","0000111111111111111111111111","0000111001101110011011100110","0000111011111110111111101111","0000111111111111111111111111","0000111011111110111111101111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110001111100011111000111","0000100000011000000110000001","0000101000011010000110100001","0000100010001000100010001000","0000011010010110100101101001","0000100011011000110110001101","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000110010101100101011001010","0000111010101110101011101010","0000101011101010111010101110","0000111111111111111111111111","0000111011101110111011101110","0000111000111110001111100011","0000111011011110110111101101","0000111110101111101011111010","0000111111101111111011111110","0000111111011111110111111101","0000111100111111001111110011","0000111110001111100011111000","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111101011111010111110101","0000111101001111010011110100","0000111110011111100111111001","0000111111111111111111111111","0000111110011111100111111001","0000110110111101101111011011","0000101100011011000110110001","0000011101010111010101110101","0000100100001001000010010000","0000100010101000101010001010","0000011101110111011101110111","0000100101111001011110010111","0000011100000111000001110000","0000010001000100010001000100","0000010001100100011001000110","0000010111000101110001011100","0000010110110101101101011011","0000010011110100111101001111","0000011101000111010001110100","0000101000101010001010100010","0000101000011010000110100001","0000100111111001111110011111","0000100010001000100010001000","0000011000000110000001100000","0000010001100100011001000110","0000001010100010101000101010","0000011001010110010101100101","0000010101010101010101010101","0000101001101010011010100110","0000011010010110100101101001","0000100000111000001110000011","0000100001101000011010000110","0000011000100110001001100010","0001000000000000000000000000","0000011001010110010101100101","0000011001000110010001100100","0000110111001101110011011100","0000011110000111100001111000","0000110000101100001011000010","0000111011011110110111101101","0000101010011010100110101001","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111001001110010011100100","0000111000101110001011100010","0000111010101110101011101010","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111011011110110111101101","0000111001111110011111100111","0000111111001111110011111100","0000111101011111010111110101","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111100011111000111110001","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111101111111011111110","0000111100101111001011110010","0000110011111100111111001111","0000010100110101001101010011","0000111001011110010111100101","0000110111101101111011011110","0000111100001111000011110000","0000110111101101111011011110","0000110011001100110011001100","0000111111111111111111111111","0000110101001101010011010100","0000111001011110010111100101","0000110101111101011111010111","0000111100001111000011110000","0000111111111111111111111111","0000111100001111000011110000","0000011100110111001101110011","0000010111100101111001011110","0000000000100000001000000010","0000000011110000111100001111","0000011010110110101101101011","0000100101001001010010010100","0000011101100111011001110110","0000100101111001011110010111","0000111001101110011011100110","0000111111111111111111111111","0000111011111110111111101111","0000111101011111010111110101","0000110110001101100011011000","0000010110110101101101011011","0000000001100000011000000110","0000010001000100010001000100","0000101001111010011110100111","0000111000111110001111100011","0000101110001011100010111000","0000101001101010011010100110","0000101111011011110110111101","0000111111101111111011111110","0000111001111110011111100111","0000110011001100110011001100","0000100001111000011110000111","0000100011111000111110001111","0000011000110110001101100011","0000110001111100011111000111","0000010000010100000101000001","0000001110010011100100111001","0000011001010110010101100101","0000010011100100111001001110","0000011010110110101101101011","0000111111101111111011111110","0000111111111111111111111111","0000111010001110100011101000","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000101001001010010010100100","0001000000000000000000000000","0000000010110000101100001011","0000101001001010010010100100","0000100110001001100010011000","0000110000011100000111000001","0000110010001100100011001000","0000111011101110111011101110","0000110011111100111111001111","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000110010111100101111001011","0000010101010101010101010101","0000100100101001001010010010","0000011110100111101001111010","0000011010000110100001101000","0000011101110111011101110111","0000111101011111010111110101","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111100111111001111110011","0000110011101100111011001110","0000111010001110100011101000","0000101100001011000010110000","0000110110001101100011011000","0000111110011111100111111001","0000111000111110001111100011","0000111011001110110011101100","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111111111111111111111111","0000111100101111001011110010","0000111010011110100111101001","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000110100111101001111010011","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000111110101111101011111010","0000111111101111111011111110","0000111101001111010011110100","0000111000011110000111100001","0000111101001111010011110100","0000111111101111111011111110","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000101111111011111110111111","0000101001111010011110100111","0000100110101001101010011010","0000100101001001010010010100","0000110000001100000011000000","0000110111101101111011011110","0000110111101101111011011110","0000101011101010111010101110","0000011010110110101101101011","0000001101100011011000110110","0000000010100000101000001010","0000000110000001100000011000","0000010110000101100001011000","0000011110000111100001111000","0000001101100011011000110110","0000010010100100101001001010","0000010110010101100101011001","0000101010001010100010101000","0000100111101001111010011110","0000011100000111000001110000","0000100001001000010010000100","0000010111100101111001011110","0000100010111000101110001011","0000000101110001011100010111","0000001100100011001000110010","0000000000110000001100000011","0000001111010011110100111101","0000010110110101101101011011","0000111000001110000011100000","0000100110111001101110011011","0000110010011100100111001001","0000110110101101101011011010","0000101110011011100110111001","0000111011111110111111101111","0000111110111111101111111011","0000111101001111010011110100","0000111010011110100111101001","0000101101011011010110110101","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000110100101101001011010010","0000101000101010001010100010","0000010111100101111001011110","0000110111101101111011011110","0000110100001101000011010000","0000111010101110101011101010","0000111111111111111111111111","0000111100101111001011110010","0000111001101110011011100110","0000111011001110110011101100","0000111010011110100111101001","0000111010101110101011101010","0000110101111101011111010111","0000111011111110111111101111","0000111110001111100011111000","0000111110101111101011111010","0000110101101101011011010110","0000011011100110111001101110","0000010011100100111001001110","0001000000000000000000000000","0000000101010001010100010101","0000100101011001010110010101","0000100011011000110110001101","0000100110101001101010011010","0000101101101011011010110110","0000111111111111111111111111","0000111110101111101011111010","0000111100001111000011110000","0000011110000111100001111000","0000001101010011010100110101","0000010000100100001001000010","0000101000001010000010100000","0000111010111110101111101011","0000111011101110111011101110","0000111100011111000111110001","0000110111001101110011011100","0000100001011000010110000101","0000011111110111111101111111","0000111111101111111011111110","0000100111001001110010011100","0000011111100111111001111110","0000100101011001010110010101","0000100010111000101110001011","0000010011110100111101001111","0000000011010000110100001101","0000001100100011001000110010","0000011010110110101101101011","0000010000110100001101000011","0000111111111111111111111111","0000111100011111000111110001","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111010001110100011101000","0000111111101111111011111110","0000000110100001101000011010","0000000000010000000100000001","0000011111110111111101111111","0000100000001000000010000000","0000011111010111110101111101","0000100000101000001010000010","0000111110001111100011111000","0000101001111010011110100111","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000110100111101001111010011","0000010001000100010001000100","0000100001011000010110000101","0000011001100110011001100110","0000011001000110010001100100","0000001100100011001000110010","0000111110101111101011111010","0000111101111111011111110111","0000111011111110111111101111","0000111111011111110111111101","0000110111001101110011011100","0000110010001100100011001000","0000111111111111111111111111","0000100100001001000010010000","0000111101001111010011110100","0000111000101110001011100010","0000111011111110111111101111","0000111110101111101011111010","0000111111011111110111111101","0000111100111111001111110011","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111101101111011011110110","0000111101011111010111110101","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111011011110110111101101","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000101110111011101110111011","0000111110101111101011111010","0000111011011110110111101101","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111001001110010011100100","0000110010011100100111001001","0000111111111111111111111111","0000111001111110011111100111","0000110110101101101011011010","0000111110011111100111111001","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111101111111011111110","0000110111011101110111011101","0000110011001100110011001100","0000101111011011110110111101","0000110011111100111111001111","0000111000001110000011100000","0000110011101100111011001110","0000101110101011101010111010","0000100111101001111010011110","0000011101000111010001110100","0000010000010100000101000001","0000011001100110011001100110","0000100000101000001010000010","0000101110101011101010111010","0000101100001011000010110000","0000100000101000001010000010","0000011001100110011001100110","0000011010000110100001101000","0000010111000101110001011100","0000011101110111011101110111","0000100010001000100010001000","0001000000000000000000000000","0001000000000000000000000000","0000010101110101011101010111","0000100011101000111010001110","0000010101010101010101010101","0000101100101011001010110010","0000101101001011010010110100","0000110000001100000011000000","0000111101001111010011110100","0000111000111110001111100011","0000111111111111111111111111","0000111111111111111111111111","0000110001001100010011000100","0000111010101110101011101010","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111100111111001111110011","0000111110011111100111111001","0000111110111111101111111011","0000111101011111010111110101","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111100001111000011110000","0000111110111111101111111011","0000111110111111101111111011","0000111100111111001111110011","0000111110001111100011111000","0000111111101111111011111110","0000111010101110101011101010","0000110010101100101011001010","0000101110001011100010111000","0000101000101010001010100010","0000011100000111000001110000","0000010110100101101001011010","0000110111111101111111011111","0000110010001100100011001000","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111010001110100011101000","0000110111111101111111011111","0000111010111110101111101011","0000111111101111111011111110","0000111110001111100011111000","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000011010100110101001101010","0000100001111000011110000111","0000000101100001011000010110","0000000111110001111100011111","0000011110100111101001111010","0000101000101010001010100010","0000100001111000011110000111","0000100110111001101110011011","0000110001011100010111000101","0000100110111001101110011011","0000011000100110001001100010","0000100000101000001010000010","0000011011000110110001101100","0000101001111010011110100111","0000100111111001111110011111","0000111111111111111111111111","0000111110011111100111111001","0000110110111101101111011011","0000110010011100100111001001","0000110001101100011011000110","0000011100000111000001110000","0000010111100101111001011110","0000011100100111001001110010","0000100101001001010010010100","0000100001001000010010000100","0000010000100100001001000010","0000001010000010100000101000","0000000011000000110000001100","0000101001111010011110100111","0000001011000010110000101100","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111111111111111111111111","0000111100111111001111110011","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000100110101001101010011010","0001000000000000000000000000","0000010101100101011001010110","0000001111010011110100111101","0000010111000101110001011100","0000001100100011001000110010","0000101100101011001010110010","0000111101001111010011110100","0000010111010101110101011101","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000110100011101000111010001","0000010100100101001001010010","0000011100110111001101110011","0000010010000100100001001000","0000011001000110010001100100","0000000010100000101000001010","0000110111101101111011011110","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000110010111100101111001011","0000111101001111010011110100","0000111111001111110011111100","0000101011101010111010101110","0000111110001111100011111000","0000110011101100111011001110","0000111110111111101111111011","0000111111101111111011111110","0000111101001111010011110100","0000111110101111101011111010","0000111111101111111011111110","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111001001110010011100100","0000111010101110101011101010","0000111010111110101111101011","0000111111111111111111111111","0000111100011111000111110001","0000111011101110111011101110","0000110111011101110111011101","0000111111111111111111111111","0000111010111110101111101011","0000110111011101110111011101","0000101011011010110110101101","0000111100011111000111110001","0000110111101101111011011110","0000111111101111111011111110","0000111111111111111111111111","0000111011111110111111101111","0000111000001110000011100000","0000101101001011010010110100","0000111111111111111111111111","0000110100011101000111010001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111011001110110011101100","0000110001111100011111000111","0000101100001011000010110000","0000011010100110101001101010","0000011100110111001101110011","0000010011110100111101001111","0000010000110100001101000011","0000011110110111101101111011","0000101010101010101010101010","0000101101001011010010110100","0000010100000101000001010000","0000001001000010010000100100","0000011000010110000101100001","0000100000001000000010000000","0000000101010001010100010101","0001000000000000000000000000","0000001100000011000000110000","0000011100110111001101110011","0000010110000101100001011000","0000010101000101010001010100","0000100010101000101010001010","0000100001001000010010000100","0000110000101100001011000010","0000111101011111010111110101","0000111101111111011111110111","0000110110001101100011011000","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111011001110110011101100","0000111100101111001011110010","0000111110011111100111111001","0000111110001111100011111000","0000111100011111000111110001","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111100111111001111110011","0000110111111101111111011111","0000110011001100110011001100","0000101111111011111110111111","0000101110101011101010111010","0000101000111010001110100011","0000101000011010000110100001","0000101011101010111010101110","0000100110001001100010011000","0000011011110110111101101111","0000011011100110111001101110","0000100011101000111010001110","0000011000110110001101100011","0001000000000000000000000000","0000001010010010100100101001","0000010101110101011101010111","0000011000010110000101100001","0000011011110110111101101111","0000010101010101010101010101","0000011111010111110101111101","0000101110101011101010111010","0000110111111101111111011111","0000111000111110001111100011","0000111110101111101011111010","0000110000111100001111000011","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111100001111000011110000","0000111010111110101111101011","0000101101111011011110110111","0000011011010110110101101101","0000011100000111000001110000","0000000010100000101000001010","0000011001010110010101100101","0000100110001001100010011000","0000001111010011110100111101","0000011101100111011001110110","0000100111011001110110011101","0000110011011100110111001101","0000101111011011110110111101","0000101110101011101010111010","0000100010001000100010001000","0000101001011010010110100101","0000111100011111000111110001","0000111101001111010011110100","0000111111101111111011111110","0000111110111111101111111011","0000110101001101010011010100","0000100100011001000110010001","0000011001010110010101100101","0000010000010100000101000001","0000011110010111100101111001","0000100001101000011010000110","0000011011000110110001101100","0000000001000000010000000100","0000000010110000101100001011","0000100011011000110110001101","0000000011100000111000001110","0000110100011101000111010001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111010101110101011101010","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111111011111110111111101","0000111100101111001011110010","0000000000010000000100000001","0000000010100000101000001010","0000000000010000000100000001","0000010011100100111001001110","0000010100000101000001010000","0000001100010011000100110001","0000101100111011001110110011","0000111001011110010111100101","0000011100100111001001110010","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111001111110011111100","0000111101011111010111110101","0000111110011111100111111001","0000110000101100001011000010","0000010111100101111001011110","0000010110010101100101011001","0000001001010010010100100101","0000010111010101110101011101","0000000010010000100100001001","0000011010100110101001101010","0000111000011110000111100001","0000111111111111111111111111","0000111100101111001011110010","0000101101101011011010110110","0000111001001110010011100100","0000110010011100100111001001","0000111001111110011111100111","0000111100011111000111110001","0000101101101011011010110110","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111111111111111111111111","0000111000111110001111100011","0000111000111110001111100011","0000111010001110100011101000","0000111110111111101111111011","0000101111001011110010111100","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000110101011101010111010101","0000111010101110101011101010","0000111111101111111011111110","0000110111101101111011011110","0000101101111011011110110111","0000110110111101101111011011","0000101110011011100110111001","0000111101111111011111110111","0000111111111111111111111111","0000111100101111001011110010","0000111100111111001111110011","0000101011101010111010101110","0000111010011110100111101001","0000101001111010011110100111","0000111110011111100111111001","0000111111111111111111111111","0000110111111101111111011111","0000111100011111000111110001","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000111100101111001011110010","0000111100001111000011110000","0000111111011111110111111101","0000111111111111111111111111","0000111101101111011011110110","0000111001111110011111100111","0000110110101101101011011010","0000110011101100111011001110","0000101001001010010010100100","0000100111111001111110011111","0000101001011010010110100101","0000101100001011000010110000","0000101100111011001110110011","0000101001001010010010100100","0000011111100111111001111110","0000000011110000111100001111","0000001111000011110000111100","0000100011111000111110001111","0000000100100001001000010010","0000000010110000101100001011","0000011010100110101001101010","0000101101101011011010110110","0000001001110010011100100111","0000010001110100011101000111","0000010001110100011101000111","0000010100000101000001010000","0000100100011001000110010001","0000100000011000000110000001","0000101001101010011010100110","0000110001011100010111000101","0000111111111111111111111111","0000110011001100110011001100","0000110101011101010111010101","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111101101111011011110110","0000111100001111000011110000","0000111010101110101011101010","0000111001101110011011100110","0000111010111110101111101011","0000111110111111101111111011","0000111001001110010011100100","0000101010011010100110101001","0000100001011000010110000101","0000011110000111100001111000","0000010100010101000101010001","0000000110110001101100011011","0000001010110010101100101011","0000011111010111110101111101","0000010110110101101101011011","0000011011000110110001101100","0000100010011000100110001001","0000101000101010001010100010","0000101010111010101110101011","0000101011101010111010101110","0000100101111001011110010111","0000011101110111011101110111","0000110010011100100111001001","0000111111111111111111111111","0000110010101100101011001010","0000111110111111101111111011","0000111011111110111111101111","0000111101111111011111110111","0000110110101101101011011010","0000110100011101000111010001","0000110000111100001111000011","0000101110101011101010111010","0000011001010110010101100101","0000001110110011101100111011","0000000011100000111000001110","0000000010100000101000001010","0000010000110100001101000011","0000100101101001011010010110","0000001111010011110100111101","0000101101001011010010110100","0000111111111111111111111111","0000110110001101100011011000","0000101111101011111010111110","0000100110001001100010011000","0000110101111101011111010111","0000111110011111100111111001","0000111110101111101011111010","0000111101101111011011110110","0000111111111111111111111111","0000111101011111010111110101","0000110101001101010011010100","0000000001010000010100000101","0000001111100011111000111110","0000001111100011111000111110","0000011111000111110001111100","0000001100110011001100110011","0000000111100001111000011110","0000001110110011101100111011","0000000011100000111000001110","0000110001011100010111000101","0000111011011110110111101101","0000111111111111111111111111","0000111111011111110111111101","0000111100001111000011110000","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111110011111100111111001","0000111111111111111111111111","0000101011101010111010101110","0000010011010100110101001101","0000001010000010100000101000","0000010011100100111001001110","0000001011000010110000101100","0000001001000010010000100100","0000010111000101110001011100","0000101100011011000110110001","0000101100111011001110110011","0000101000101010001010100010","0000111011101110111011101110","0000111100011111000111110001","0000111011101110111011101110","0000111111111111111111111111","0000111110101111101011111010","0000101011101010111010101110","0000001011010010110100101101","0000010110010101100101011001","0000010001110100011101000111","0000011110010111100101111001","0000010011100100111001001110","0000010100100101001001010010","0000100100101001001010010010","0000101011111010111110101111","0000110110011101100111011001","0000110100101101001011010010","0000110100101101001011010010","0000110100101101001011010010","0000110011101100111011001110","0000110011111100111111001111","0000101101111011011110110111","0000111001001110010011100100","0000111011011110110111101101","0000111111111111111111111111","0000111101011111010111110101","0000110110001101100011011000","0000111110001111100011111000","0000111111011111110111111101","0000111100111111001111110011","0000110010101100101011001010","0000111000001110000011100000","0000110111011101110111011101","0000110100001101000011010000","0000110010001100100011001000","0000111100111111001111110011","0000111101111111011111110111","0000110111111101111111011111","0000110111011101110111011101","0000111110101111101011111010","0000101111101011111010111110","0000101101111011011110110111","0000101111111011111110111111","0000110010101100101011001010","0000111111111111111111111111","0000110110001101100011011000","0000111111111111111111111111","0000101001011010010110100101","0000111001111110011111100111","0000101010011010100110101001","0000111111111111111111111111","0000111111111111111111111111","0000101111001011110010111100","0000111111101111111011111110","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111011101110111011101110","0000111111001111110011111100","0000111111111111111111111111","0000111010101110101011101010","0000101100001011000010110000","0000101101111011011110110111","0000110100011101000111010001","0000111001001110010011100100","0000111011101110111011101110","0000110101111101011111010111","0000100111111001111110011111","0000110011001100110011001100","0000111000101110001011100010","0000110010011100100111001001","0000011111010111110101111101","0000000100100001001000010010","0000001110000011100000111000","0000011001110110011101100111","0000001000010010000100100001","0000000011110000111100001111","0000001110110011101100111011","0000010001100100011001000110","0000010011010100110101001101","0000001100010011000100110001","0000001101010011010100110101","0000001000100010001000100010","0000001000110010001100100011","0000011101010111010101110101","0000010101100101011001010110","0000100100101001001010010010","0000100110111001101110011011","0000100101101001011010010110","0000110001011100010111000101","0000111101101111011011110110","0000111111111111111111111111","0000111110111111101111111011","0000111100011111000111110001","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000101101001011010010110100","0000101001101010011010100110","0000010100100101001001010010","0000000010010000100100001001","0000001111110011111100111111","0000011100000111000001110000","0000011010110110101101101011","0000101000101010001010100010","0000100011011000110110001101","0000100001101000011010000110","0000100001101000011010000110","0000100001001000010010000100","0000100100011001000110010001","0000100111011001110110011101","0000100110011001100110011001","0000110100101101001011010010","0000111001011110010111100101","0000100011101000111010001110","0000110011011100110111001101","0000101100011011000110110001","0000111100001111000011110000","0000110010001100100011001000","0000111101101111011011110110","0000111110101111101011111010","0000111100101111001011110010","0000110101101101011011010110","0000101000001010000010100000","0000101011001010110010101100","0000000101000001010000010100","0000000011100000111000001110","0000000000100000001000000010","0000001110000011100000111000","0000110110011101100111011001","0000011101010111010101110101","0000110110001101100011011000","0000111111001111110011111100","0000110011111100111111001111","0000110010111100101111001011","0000100111001001110010011100","0000110101111101011111010111","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000101100111011001110110011","0000010111100101111001011110","0000001001000010010000100100","0000001001110010011100100111","0000011110100111101001111010","0000000111010001110100011101","0000101000001010000010100000","0000000011010000110100001101","0000101110011011100110111001","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111100011111000111110001","0000111100001111000011110000","0000011011010110110101101101","0000001000100010001000100010","0000010101100101011001010110","0000000000100000001000000010","0000000001100000011000000110","0000000110100001101000011010","0000010101000101010001010100","0000011011100110111001101110","0000101000111010001110100011","0000100010101000101010001010","0000110011001100110011001100","0000111011111110111111101111","0000111000111110001111100011","0000110010101100101011001010","0000100010011000100110001001","0000110010001100100011001000","0000001010110010101100101011","0000010000110100001101000011","0000011100010111000101110001","0000001100000011000000110000","0000001000000010000000100000","0000011111100111111001111110","0000011101110111011101110111","0000100111011001110110011101","0000100001011000010110000101","0000101011111010111110101111","0000101100101011001010110010","0000110011111100111111001111","0000101001101010011010100110","0000101010011010100110101001","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000101111111011111110111111","0000111111001111110011111100","0000111111101111111011111110","0000111110101111101011111010","0000111000001110000011100000","0000110000101100001011000010","0000101001101010011010100110","0000011110110111101101111011","0000011101110111011101110111","0000011101110111011101110111","0000011010010110100101101001","0000100011101000111010001110","0000011100100111001001110010","0000110011101100111011001110","0000101110001011100010111000","0000101010011010100110101001","0000100010101000101010001010","0000110001011100010111000101","0000111111111111111111111111","0000101101101011011010110110","0000111100011111000111110001","0000101101101011011010110110","0000111011001110110011101100","0000101010101010101010101010","0000111111111111111111111111","0000111101111111011111110111","0000101101001011010010110100","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111001011110010111100101","0000111000001110000011100000","0000110100111101001111010011","0000110001011100010111000101","0000100010011000100110001001","0000100010111000101110001011","0000100110111001101110011011","0000110001111100011111000111","0000110111001101110011011100","0000110110001101100011011000","0000110110001101100011011000","0000110001001100010011000100","0000111011011110110111101101","0000101000011010000110100001","0001000000000000000000000000","0000001010110010101100101011","0000010000110100001101000011","0001000000000000000000000000","0001000000000000000000000000","0000000101100001011000010110","0000000100100001001000010010","0000001000100010001000100010","0000011110010111100101111001","0000001000110010001100100011","0000000100000001000000010000","0000010101100101011001010110","0000010001110100011101000111","0000011000110110001101100011","0000011010000110100001101000","0000010011110100111101001111","0000011111010111110101111101","0000101001111010011110100111","0000110011011100110111001101","0000110111011101110111011101","0000111011001110110011101100","0000111110111111101111111011","0000111100101111001011110010","0000110110111101101111011011","0000110101101101011011010110","0000110010101100101011001010","0000110111101101111011011110","0000110101111101011111010111","0000110000011100000111000001","0000101010101010101010101010","0000011110000111100001111000","0000010111000101110001011100","0000010100010101000101010001","0000000101010001010100010101","0001000000000000000000000000","0000010010010100100101001001","0000110001101100011011000110","0000111010011110100111101001","0000110010001100100011001000","0000101100101011001010110010","0000100001111000011110000111","0000101001101010011010100110","0000110011111100111111001111","0000111010101110101011101010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000110111011101110111011101","0000110101101101011011010110","0000101111111011111110111111","0000011011110110111101101111","0000101101111011011110110111","0000111011101110111011101110","0000101010101010101010101010","0000111101101111011011110110","0000111010001110100011101000","0000111111111111111111111111","0000111111001111110011111100","0000110110111101101111011011","0000110011011100110111001101","0000000110100001101000011010","0001000000000000000000000000","0000011111110111111101111111","0000001000010010000100100001","0000100111001001110010011100","0000101111111011111110111111","0000110000001100000011000000","0000111011111110111111101111","0000110000101100001011000010","0000110011101100111011001110","0000101111011011110110111101","0000111100111111001111110011","0000110101011101010111010101","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000101010011010100110101001","0000010101010101010101010101","0001000000000000000000000000","0000001101110011011100110111","0000010000010100000101000001","0000100010101000101010001010","0000100000101000001010000010","0000100111001001110010011100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000110000001100000011000000","0000001100100011001000110010","0000001011000010110000101100","0000010011010100110101001101","0000011000110110001101100011","0000000100000001000000010000","0001000000000000000000000000","0000001100100011001000110010","0000010011100100111001001110","0000100010001000100010001000","0000011111110111111101111111","0000101001101010011010100110","0000101010111010101110101011","0000101011001010110010101100","0000100011101000111010001110","0000101110111011101110111011","0000010001010100010101000101","0000010111100101111001011110","0000001100000011000000110000","0000011000110110001101100011","0000000011100000111000001110","0000010111000101110001011100","0000011100010111000101110001","0000011100000111000001110000","0000010111100101111001011110","0000100000101000001010000010","0000100010101000101010001010","0000100100001001000010010000","0000101110101011101010111010","0000101101011011010110110101","0000111101011111010111110101","0000110101001101010011010100","0000111111111111111111111111","0000111000011110000111100001","0000110111111101111111011111","0000101001011010010110100101","0000111100101111001011110010","0000111011001110110011101100","0000111111111111111111111111","0000110010001100100011001000","0000100010001000100010001000","0000011110100111101001111010","0000010000010100000101000001","0000011001000110010001100100","0000100000111000001110000011","0000101100001011000010110000","0000011000010110000101100001","0000011001000110010001100100","0000100000011000000110000001","0000011011100110111001101110","0000010110000101100001011000","0000011011010110110101101101","0000111111111111111111111111","0000101000011010000110100001","0000101110001011100010111000","0000100100101001001010010010","0000110101001101010011010100","0000110110011101100111011001","0000111011101110111011101110","0000111011111110111111101111","0000101101111011011110110111","0000111110101111101011111010","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111101001111010011110100","0000111111011111110111111101","0000111100001111000011110000","0000111011011110110111101101","0000111101011111010111110101","0000111011001110110011101100","0000110110101101101011011010","0000101100011011000110110001","0000110011111100111111001111","0000101010011010100110101001","0000011110110111101101111011","0000101000011010000110100001","0000101100101011001010110010","0000101110101011101010111010","0000110110101101101011011010","0000110111001101110011011100","0000110000111100001111000011","0000100011011000110110001101","0000001100110011001100110011","0000000010000000100000001000","0000010100110101001101010011","0000001000010010000100100001","0000001100010011000100110001","0000001101110011011100110111","0000011001100110011001100110","0000010010010100100101001001","0000000011110000111100001111","0000000010000000100000001000","0000000100100001001000010010","0000001111110011111100111111","0000010001010100010101000101","0000010101110101011101010111","0000001010110010101100101011","0000010100100101001001010010","0000001000100010001000100010","0000001011010010110100101101","0000010000010100000101000001","0000010011000100110001001100","0000001111000011110000111100","0000001000000010000000100000","0000000101000001010000010100","0000000110100001101000011010","0000000001000000010000000100","0000001001000010010000100100","0000000110110001101100011011","0000000111010001110100011101","0000000101010001010100010101","0000000101000001010000010100","0000010011010100110101001101","0000011010010110100101101001","0000011010100110101001101010","0000001111100011111000111110","0000101101101011011010110110","0000111110011111100111111001","0000110110011101100111011001","0000111010101110101011101010","0000111001101110011011100110","0000110010101100101011001010","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111110101111101011111010","0000111110001111100011111000","0000111101111111011111110111","0000111110001111100011111000","0000111011101110111011101110","0000110101011101010111010101","0000010000110100001101000011","0000110101011101010111010101","0000100100011001000110010001","0000111111111111111111111111","0000111001011110010111100101","0000110010101100101011001010","0000110101111101011111010111","0000110011001100110011001100","0000111001111110011111100111","0000110001001100010011000100","0000010011000100110001001100","0000000010000000100000001000","0000011100100111001001110010","0000100010011000100110001001","0000000111110001111100011111","0000100010111000101110001011","0000100011001000110010001100","0000110000101100001011000010","0000101111011011110110111101","0000101110111011101110111011","0000110010001100100011001000","0000110001011100010111000101","0000110101101101011011010110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000110001001100010011000100","0000110011011100110111001101","0000010101100101011001010110","0000001011100010111000101110","0000010101100101011001010110","0000001001010010010100100101","0000101011001010110010101100","0000001101100011011000110110","0000111101111111011111110111","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000011111000111110001111100","0001000000000000000000000000","0000100110001001100010011000","0000100100111001001110010011","0000101101001011010010110100","0000011001100110011001100110","0001000000000000000000000000","0000001010000010100000101000","0000001110010011100100111001","0000010100000101000001010000","0000010011110100111101001111","0000011011100110111001101110","0000011100000111000001110000","0000110100001101000011010000","0000100010111000101110001011","0000101001101010011010100110","0000010111100101111001011110","0000011111000111110001111100","0000010000110100001101000011","0000010110110101101101011011","0000001001110010011100100111","0000100111101001111010011110","0000100110111001101110011011","0000001100010011000100110001","0000010011100100111001001110","0000100001101000011010000110","0000011110000111100001111000","0000100111101001111010011110","0000110010111100101111001011","0000111010111110101111101011","0000111100111111001111110011","0000101110011011100110111001","0000111000111110001111100011","0000111011111110111111101111","0000110111101101111011011110","0000100110101001101010011010","0000101100001011000010110000","0000111000101110001011100010","0000111111001111110011111100","0000111111111111111111111111","0000101100101011001010110010","0000100011011000110110001101","0000000111000001110000011100","0000001011000010110000101100","0000001011110010111100101111","0000000101010001010100010101","0000000100000001000000010000","0000001101010011010100110101","0000001101000011010000110100","0000000111000001110000011100","0000001100010011000100110001","0000110010001100100011001000","0000100111111001111110011111","0000101010011010100110101001","0000011101010111010101110101","0000011110010111100101111001","0000110010011100100111001001","0000111011011110110111101101","0000111101111111011111110111","0000110010001100100011001000","0000111111001111110011111100","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111001111110011111100111","0000110101101101011011010110","0000110111011101110111011101","0000111111111111111111111111","0000110001001100010011000100","0000110011011100110111001101","0000110111011101110111011101","0000001110010011100100111001","0000100111101001111010011110","0000100100101001001010010010","0000111101101111011011110110","0000111111111111111111111111","0000101001001010010010100100","0000100011001000110010001100","0000011000110110001101100011","0001000000000000000000000000","0000010110010101100101011001","0000001011000010110000101100","0000001010000010100000101000","0000010011100100111001001110","0000011111110111111101111111","0000001110100011101000111010","0000100000011000000110000001","0000011000000110000001100000","0000011110000111100001111000","0000010010100100101001001010","0000010110100101101001011010","0000001100010011000100110001","0000000111000001110000011100","0001000000000000000000000000","0001000000000000000000000000","0000001111010011110100111101","0000010111000101110001011100","0000001101000011010000110100","0000000100100001001000010010","0000001100010011000100110001","0000011011110110111101101111","0000100101111001011110010111","0000100110011001100110011001","0000101010101010101010101010","0000100111001001110010011100","0000100000101000001010000010","0000101110001011100010111000","0000101100111011001110110011","0000011011010110110101101101","0000100100111001001110010011","0000101100001011000010110000","0000111000111110001111100011","0000110101101101011011010110","0000111000001110000011100000","0000111110001111100011111000","0000111100111111001111110011","0000111110101111101011111010","0000111100001111000011110000","0000111110101111101011111010","0000111110101111101011111010","0000111100001111000011110000","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110001111100011111000111","0000010001110100011101000111","0000101001101010011010100110","0000100110111001101110011011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000001110000011100000","0000110111101101111011011110","0000110000001100000011000000","0000100101001001010010010100","0000000100000001000000010000","0000000001010000010100000101","0000001011000010110000101100","0000011001010110010101100101","0000011010100110101001101010","0000001110100011101000111010","0000101001101010011010100110","0000110110011101100111011001","0000110010101100101011001010","0000100110011001100110011001","0000110011111100111111001111","0000101011111010111110101111","0000111110101111101011111010","0000111110001111100011111000","0000111101111111011111110111","0000111111111111111111111111","0000101111011011110110111101","0000110010111100101111001011","0000010110000101100001011000","0000011000010110000101100001","0000000111010001110100011101","0000011110010111100101111001","0000010111000101110001011100","0000100010011000100110001001","0000111101111111011111110111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000110110011101100111011001","0000000111110001111100011111","0000001011010010110100101101","0000110101111101011111010111","0000101111101011111010111110","0000111001001110010011100100","0000100110011001100110011001","0000000010110000101100001011","0000000001000000010000000100","0000001010000010100000101000","0000010010010100100101001001","0000100011101000111010001110","0000101100001011000010110000","0000100011001000110010001100","0000111010001110100011101000","0000110000111100001111000011","0000011100000111000001110000","0000100101101001011010010110","0000010101000101010001010100","0000010111000101110001011100","0000001100010011000100110001","0000011111000111110001111100","0000100110101001101010011010","0000011001110110011101100111","0000011101010111010101110101","0000011111100111111001111110","0000010000010100000101000001","0000011000010110000101100001","0000101110011011100110111001","0000100011101000111010001110","0000111010101110101011101010","0000111001011110010111100101","0000101000111010001110100011","0000101111111011111110111111","0000110000001100000011000000","0000101011101010111010101110","0000110001001100010011000100","0000100010111000101110001011","0000100000011000000110000001","0000100100011001000110010001","0000010011000100110001001100","0001000000000000000000000000","0000000000110000001100000011","0000000001010000010100000101","0000000011110000111100001111","0000001101100011011000110110","0000010101000101010001010100","0000000100000001000000010000","0000001010010010100100101001","0000000000010000000100000001","0000000110000001100000011000","0000010110100101101001011010","0000101100011011000110110001","0000100111011001110110011101","0000011001010110010101100101","0000010001100100011001000110","0000100010111000101110001011","0000110100011101000111010001","0000111111111111111111111111","0000110100001101000011010000","0000111100111111001111110011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111100001111000011110000","0000111010011110100111101001","0000111111111111111111111111","0000110001001100010011000100","0000101000101010001010100010","0000100110011001100110011001","0000010011100100111001001110","0000011111010111110101111101","0000111100001111000011110000","0000111110011111100111111001","0000110010011100100111001001","0000100011001000110010001100","0000010101010101010101010101","0000000110100001101000011010","0000010101100101011001010110","0000000111110001111100011111","0000000010000000100000001000","0000011001010110010101100101","0000011110000111100001111000","0000010011110100111101001111","0000010111000101110001011100","0000010000010100000101000001","0000010111000101110001011100","0000011010100110101001101010","0000101010011010100110101001","0000011010100110101001101010","0000101110101011101010111010","0000111111111111111111111111","0000110101001101010011010100","0000110000001100000011000000","0000101110111011101110111011","0000110010011100100111001001","0000110010101100101011001010","0000101100001011000010110000","0000100100101001001010010010","0000100000111000001110000011","0000100000101000001010000010","0000011110010111100101111001","0000100011101000111010001110","0000101001001010010010100100","0000011011010110110101101101","0000011111100111111001111110","0000110111101101111011011110","0000110011111100111111001111","0000101101101011011010110110","0000101110101011101010111010","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111100101111001011110010","0000111101101111011011110110","0000111111111111111111111111","0000110101101101011011010110","0000100001011000010110000101","0000011100010111000101110001","0000001110100011101000111010","0000110110001101100011011000","0000111101011111010111110101","0000111100101111001011110010","0000111110101111101011111010","0000111011101110111011101110","0000101010011010100110101001","0000101110001011100010111000","0000011010100110101001101010","0000000101100001011000010110","0001000000000000000000000000","0000000110000001100000011000","0000010100010101000101010001","0000011101100111011001110110","0000011110000111100001111000","0000010011000100110001001100","0000110001111100011111000111","0000110011011100110111001101","0000101101011011010110110101","0000101100101011001010110010","0000111011111110111111101111","0000111111011111110111111101","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000110111101101111011011110","0000100110011001100110011001","0000010101000101010001010100","0000011100100111001001110010","0000001010010010100100101001","0000101000011010000110100001","0000010010010100100101001001","0000110110011101100111011001","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111101001111010011110100","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000101001111010011110100111","0001000000000000000000000000","0000100001011000010110000101","0000111111111111111111111111","0000110010011100100111001001","0000110101011101010111010101","0000110010111100101111001011","0000011110100111101001111010","0000001001000010010000100100","0000000111100001111000011110","0000000010110000101100001011","0000010101110101011101010111","0000110101101101011011010110","0000110111111101111111011111","0000110001011100010111000101","0000100011111000111110001111","0000011000000110000001100000","0000101000111010001110100011","0000010010000100100001001000","0000001011110010111100101111","0000011001000110010001100100","0000110100101101001011010010","0000100000001000000010000000","0000100000111000001110000011","0000100001001000010010000100","0000011011100110111001101110","0001000000000000000000000000","0000001111010011110100111101","0000100000001000000010000000","0000110111101101111011011110","0000110100111101001111010011","0000110110101101101011011010","0000101000011010000110100001","0000011110010111100101111001","0000100010101000101010001010","0000011110110111101101111011","0000100000011000000110000001","0000010100110101001101010011","0001000000000000000000000000","0000010010000100100001001000","0000010111110101111101011111","0000101100101011001010110010","0000100111111001111110011111","0000010100110101001101010011","0000011000110110001101100011","0000100010001000100010001000","0000011101010111010101110101","0000100010001000100010001000","0000010100100101001001010010","0001000000000000000000000000","0000001010110010101100101011","0000010011100100111001001110","0000100000111000001110000011","0000011101010111010101110101","0000000110010001100100011001","0000100101001001010010010100","0000100000011000000110000001","0000111111101111111011111110","0000110001101100011011000110","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111100011111000111110001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000110101111101011111010111","0000111000011110000111100001","0000100100001001000010010000","0000010110100101101001011010","0000110110111101101111011011","0000111001101110011011100110","0000111000111110001111100011","0000101111101011111010111110","0000110000111100001111000011","0000100100001001000010010000","0000001101100011011000110110","0000011101100111011001110110","0000001010100010101000101010","0001000000000000000000000000","0000000101000001010000010100","0000011001110110011101100111","0000001111000011110000111100","0000001010110010101100101011","0000001111000011110000111100","0000001010110010101100101011","0000010100110101001101010011","0000010001110100011101000111","0000011001000110010001100100","0000101110001011100010111000","0000110000101100001011000010","0000110010001100100011001000","0000111000011110000111100001","0000111000111110001111100011","0000110010101100101011001010","0000110000011100000111000001","0000110010111100101111001011","0000110000101100001011000010","0000101001111010011110100111","0000100110111001101110011011","0000100010011000100110001001","0000100101101001011010010110","0000100000111000001110000011","0000100000001000000010000000","0000100111111001111110011111","0000101011101010111010101110","0000110011101100111011001110","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111001111110011111100111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111111001111110011111100","0000111010111110101111101011","0000111011011110110111101101","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000100000101000001010000010","0000100010101000101010001010","0000001110100011101000111010","0000011001010110010101100101","0000111110011111100111111001","0000111010001110100011101000","0000111001011110010111100101","0000110111001101110011011100","0000111000011110000111100001","0000111111111111111111111111","0000101010011010100110101001","0000011011110110111101101111","0001000000000000000000000000","0000010101110101011101010111","0000001100000011000000110000","0000010001010100010101000101","0000011101010111010101110101","0000100100101001001010010010","0000100000011000000110000001","0000011001010110010101100101","0000011101110111011101110111","0000101001011010010110100101","0000100111101001111010011110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000111001111110011111100111","0000101001101010011010100110","0000011011010110110101101101","0000100100011001000110010001","0000011010110110101101101011","0000100100001001000010010000","0000010011010100110101001101","0000111110011111100111111001","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111110011111100111111001","0000111111111111111111111111","0000010101000101010001010100","0000011001110110011101100111","0000101001101010011010100110","0000111101111111011111110111","0000111101011111010111110101","0000111000001110000011100000","0000110101001101010011010100","0000101000101010001010100010","0000101001011010010110100101","0000011111110111111101111111","0000000111010001110100011101","0000000100110001001100010011","0000000001000000010000000100","0000001000010010000100100001","0000001011110010111100101111","0000001111010011110100111101","0000000011110000111100001111","0000100101111001011110010111","0000001011010010110100101101","0000000001110000011100000111","0000100001101000011010000110","0000011000100110001001100010","0000011010000110100001101000","0000001100010011000100110001","0000011111000111110001111100","0000010010110100101101001011","0000001110100011101000111010","0000011010000110100001101000","0000011111010111110101111101","0000111010011110100111101001","0000110000001100000011000000","0000101000001010000010100000","0000101000011010000110100001","0000011010000110100001101000","0000001111010011110100111101","0000001001110010011100100111","0000001101010011010100110101","0000010000010100000101000001","0000010101000101010001010100","0000100000001000000010000000","0000100011001000110010001100","0000110010001100100011001000","0000101011111010111110101111","0000100101001001010010010100","0000100010001000100010001000","0000101111111011111110111111","0000101111001011110010111100","0000101111111011111110111111","0000011000100110001001100010","0000000001000000010000000100","0000001000110010001100100011","0000010001110100011101000111","0000011010100110101001101010","0000010001010100010101000101","0000010011110100111101001111","0000010111100101111001011110","0000110001011100010111000101","0000101110101011101010111010","0000111010011110100111101001","0000111101001111010011110100","0000111111101111111011111110","0000111101001111010011110100","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000101100001011000010110000","0000110010101100101011001010","0000110100001101000011010000","0000111000001110000011100000","0000101000101010001010100010","0000100010101000101010001010","0000101010101010101010101010","0000110000001100000011000000","0000101001111010011110100111","0000101100001011000010110000","0000100111001001110010011100","0000101011001010110010101100","0000010010010100100101001001","0000011101000111010001110100","0000010001000100010001000100","0000000001010000010100000101","0000000100000001000000010000","0000101101111011011110110111","0000011010000110100001101000","0000000111100001111000011110","0000010011100100111001001110","0000001101010011010100110101","0000100010111000101110001011","0000010110100101101001011010","0000010010100100101001001010","0000011111000111110001111100","0000110101101101011011010110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000110011101100111011001110","0000101010011010100110101001","0000100101011001010110010101","0000100100011001000110010001","0000100001101000011010000110","0000100101101001011010010110","0000100100101001001010010010","0000101101001011010010110100","0000110111101101111011011110","0000111011101110111011101110","0000111111111111111111111111","0000111111101111111011111110","0000111011011110110111101101","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111110101111101011111010","0000111111111111111111111111","0000111011101110111011101110","0000101010011010100110101001","0000100111011001110110011101","0000010011010100110101001101","0000001100010011000100110001","0000111110101111101011111010","0000110001101100011011000110","0000111011011110110111101101","0000111101011111010111110101","0000110101111101011111010111","0000101111011011110110111101","0000101101011011010110110101","0000011000010110000101100001","0000001001010010010100100101","0000010000000100000001000000","0000100111111001111110011111","0000010110000101100001011000","0000000000010000000100000001","0001000000000000000000000000","0000011001110110011101100111","0000011010000110100001101000","0000101011111010111110101111","0000101110011011100110111001","0000100111101001111010011110","0000110111011101110111011101","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000111000001110000011100000","0000101100001011000010110000","0000101010101010101010101010","0000100001001000010010000100","0000100001101000011010000110","0000001111010011110100111101","0000101011101010111010101110","0000111101001111010011110100","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111110001111100011111000","0000111111111111111111111111","0000110010001100100011001000","0000000111100001111000011110","0000101000111010001110100011","0000111000001110000011100000","0000111110001111100011111000","0000111001011110010111100101","0000110110011101100111011001","0000101101001011010010110100","0000100110101001101010011010","0000011111100111111001111110","0000101000011010000110100001","0000110100011101000111010001","0000101001011010010110100101","0000011101100111011001110110","0000011001010110010101100101","0000011011010110110101101101","0000010110000101100001011000","0000011010010110100101101001","0000010101110101011101010111","0000001000110010001100100011","0000000101000001010000010100","0000101001101010011010100110","0000011110110111101101111011","0000011110100111101001111010","0000011010010110100101101001","0000011111010111110101111101","0000011011100110111001101110","0000010000110100001101000011","0000001111100011111000111110","0000010011100100111001001110","0000011110110111101101111011","0000010010000100100001001000","0000000110010001100100011001","0000001111100011111000111110","0000010110110101101101011011","0000100011101000111010001110","0000101110001011100010111000","0000110100101101001011010010","0000101011111010111110101111","0000101100011011000110110001","0000111000101110001011100010","0000111100001111000011110000","0000111111111111111111111111","0000100111101001111010011110","0000101000101010001010100010","0000110011011100110111001101","0000110000011100000111000001","0000111101101111011011110110","0000101111001011110010111100","0000100010111000101110001011","0000000100110001001100010011","0000001000010010000100100001","0000010100110101001101010011","0000010011100100111001001110","0000011011100110111001101110","0000000101000001010000010100","0000100010011000100110001001","0000101101101011011010110110","0000111101011111010111110101","0000111000111110001111100011","0000111001111110011111100111","0000111110001111100011111000","0000111111111111111111111111","0000111100101111001011110010","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111000101110001011100010","0000110110101101101011011010","0000111101101111011011110110","0000111101001111010011110100","0000111011111110111111101111","0000110100001101000011010000","0000101011011010110110101101","0000100011011000110110001101","0000101101011011010110110101","0000010001000100010001000100","0000101011111010111110101111","0000101001101010011010100110","0000100001001000010010000100","0000100110011001100110011001","0000100111011001110110011101","0000010101100101011001010110","0000010010000100100001001000","0000000000010000000100000001","0000010110000101100001011000","0000111000101110001011100010","0000100001001000010010000100","0000011001010110010101100101","0000011100100111001001110010","0000100010001000100010001000","0000101000101010001010100010","0000010011100100111001001110","0000100101011001010110010101","0000111001011110010111100101","0000100110101001101010011010","0000110111111101111111011111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111101111111011111110111","0000111100111111001111110011","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111101111111011111110","0000111010101110101011101010","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111010001110100011101000","0000110000101100001011000010","0000111011101110111011101110","0000111111101111111011111110","0000101101011011010110110101","0000100101011001010110010101","0000011010000110100001101000","0000000101010001010100010101","0000101110001011100010111000","0000110101011101010111010101","0000110011001100110011001100","0000111011001110110011101100","0000111111101111111011111110","0000111101011111010111110101","0000111011111110111111101111","0000100100001001000010010000","0000010110100101101001011010","0000000000110000001100000011","0000010101100101011001010110","0000011000100110001001100010","0000011101100111011001110110","0000001010010010100100101001","0000000010110000101100001011","0000010010110100101101001011","0000000111100001111000011110","0000010101110101011101010111","0000100000111000001110000011","0000101100111011001110110011","0000110110011101100111011001","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111011101110111011101110","0000111101101111011011110110","0000111011101110111011101110","0000011100110111001101110011","0000110111101101111011011110","0000100110111001101110011011","0000011101010111010101110101","0000001001100010011000100110","0000111001001110010011100100","0000111111111111111111111111","0000111111001111110011111100","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000011011010110110101101101","0000011011010110110101101101","0000111001111110011111100111","0000111001001110010011100100","0000110111001101110011011100","0000101111001011110010111100","0000011010110110101101101011","0000100000011000000110000001","0000100000011000000110000001","0000101100101011001010110010","0000110101001101010011010100","0000111100001111000011110000","0000111111111111111111111111","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000111111011111110111111101","0000111010101110101011101010","0000111100001111000011110000","0000101100001011000010110000","0000011101000111010001110100","0000100111001001110010011100","0000101000001010000010100000","0000100000111000001110000011","0000100110111001101110011011","0000100000011000000110000001","0000100010011000100110001001","0000011100100111001001110010","0000010010000100100001001000","0000011010010110100101101001","0000011100000111000001110000","0000101010111010101110101011","0000110111011101110111011101","0000111001111110011111100111","0000110010111100101111001011","0000110010011100100111001001","0000100011101000111010001110","0000100111111001111110011111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111010001110100011101000","0000110111111101111111011111","0000100110111001101110011011","0000110101111101011111010111","0000101010111010101110101011","0000111110011111100111111001","0000111001011110010111100101","0000110010011100100111001001","0000101101101011011010110110","0000001011000010110000101100","0000000100000001000000010000","0000010011100100111001001110","0000011100010111000101110001","0000001110000011100000111000","0000010110110101101101011011","0000100100111001001110010011","0000101110111011101110111011","0000111110001111100011111000","0000101111101011111010111110","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000110110011101100111011001","0000010101110101011101010111","0000011110110111101101111011","0000100010111000101110001011","0000100100011001000110010001","0000010110100101101001011010","0000101111001011110010111100","0000101101101011011010110110","0000100000011000000110000001","0000101001111010011110100111","0000010101110101011101010111","0000001101110011011100110111","0001000000000000000000000000","0000010100000101000001010000","0000111010101110101011101010","0000011111000111110001111100","0000101101001011010010110100","0000100110111001101110011011","0000011100100111001001110010","0000101101011011010110110101","0000110010011100100111001001","0000110101101101011011010110","0000111011101110111011101110","0000110111101101111011011110","0000100110111001101110011011","0000110011101100111011001110","0000111110011111100111111001","0000111111101111111011111110","0000111110001111100011111000","0000111111001111110011111100","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111100001111000011110000","0000111011101110111011101110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111011101110111011101110","0000111111011111110111111101","0000111111101111111011111110","0000111111001111110011111100","0000111111111111111111111111","0000111111001111110011111100","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101100011011000110110001","0000111010001110100011101000","0000111111111111111111111111","0000101001111010011110100111","0000101110001011100010111000","0000100011101000111010001110","0000000001010000010100000101","0000100000011000000110000001","0000110001111100011111000111","0000101010111010101110101011","0000110010011100100111001001","0000110110001101100011011000","0000111111101111111011111110","0000110110011101100111011001","0000101011111010111110101111","0000011111110111111101111111","0000000001010000010100000101","0000000101000001010000010100","0000010100100101001001010010","0000011011000110110001101100","0000100000111000001110000011","0000100001011000010110000101","0000001110000011100000111000","0000001000110010001100100011","0000010101110101011101010111","0000000110110001101100011011","0000001010100010101000101010","0000010010000100100001001000","0000011111100111111001111110","0000111010001110100011101000","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111100001111000011110000","0000101101011011010110110101","0000100110001001100010011000","0000101101011011010110110101","0000110000001100000011000000","0000000111010001110100011101","0000011110110111101101111011","0000111100111111001111110011","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000110110101101101011011010","0000000100100001001000010010","0000110101101101011011010110","0000110110011101100111011001","0000110000001100000011000000","0000010111110101111101011111","0000011100100111001001110010","0000100001001000010010000100","0000110100001101000011010000","0000111010111110101111101011","0000111011011110110111101101","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000111111101111111011111110","0000111111101111111011111110","0000111111001111110011111100","0000111011111110111111101111","0000111111011111110111111101","0000111010101110101011101010","0000100111111001111110011111","0000100000111000001110000011","0000100111101001111010011110","0000111001001110010011100100","0000100010001000100010001000","0000100111011001110110011101","0000100101011001010110010101","0000100000111000001110000011","0000101010011010100110101001","0000100110011001100110011001","0000100001111000011110000111","0000011111000111110001111100","0000011111100111111001111110","0000101000001010000010100000","0000100111111001111110011111","0000110101001101010011010100","0000110111001101110011011100","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000110110111101101111011011","0000110110001101100011011000","0000111000001110000011100000","0000110111101101111011011110","0000111110111111101111111011","0000110000011100000111000001","0000111111011111110111111101","0000110001001100010011000100","0000010100010101000101010001","0000000001010000010100000101","0000011001100110011001100110","0000011010000110100001101000","0000010001110100011101000111","0000010100000101000001010000","0000100110011001100110011001","0000111010001110100011101000","0000110100101101001011010010","0000110001001100010011000100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111010001110100011101000","0000111001001110010011100100","0000111011101110111011101110","0000110010011100100111001001","0000100000111000001110000011","0000001110100011101000111010","0000011000100110001001100010","0000101001111010011110100111","0000011111100111111001111110","0000101010011010100110101001","0000110110011101100111011001","0000011101100111011001110110","0000100000101000001010000010","0000010000110100001101000011","0000001110010011100100111001","0000000101110001011100010111","0000010011110100111101001111","0000100010011000100110001001","0000011010000110100001101000","0000101001101010011010100110","0000101001101010011010100110","0000110100101101001011010010","0000111110011111100111111001","0000111110101111101011111010","0000111110011111100111111001","0000111110101111101011111010","0000110101111101011111010111","0000110111111101111111011111","0000110011011100110111001101","0000110100111101001111010011","0000111100111111001111110011","0000111111111111111111111111","0000111101011111010111110101","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100001111000011110000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100111111001111110011","0000111100101111001011110010","0000111111101111111011111110","0000111101111111011111110111","0000110111101101111011011110","0000111101011111010111110101","0000111010011110100111101001","0000100111011001110110011101","0000110100101101001011010010","0000101011011010110110101101","0000000011010000110100001101","0000010111010101110101011101","0000101111001011110010111100","0000101100101011001010110010","0000101011101010111010101110","0000110000001100000011000000","0000111100111111001111110011","0000110111101101111011011110","0000011100000111000001110000","0000011010000110100001101000","0000010000000100000001000000","0000000101010001010100010101","0000010110100101101001011010","0000100001001000010010000100","0000100001111000011110000111","0000011100100111001001110010","0000100010101000101010001010","0000101100001011000010110000","0000011001100110011001100110","0000000001010000010100000101","0000001100110011001100110011","0000000110100001101000011010","0000001001100010011000100110","0000010110110101101101011011","0000100111111001111110011111","0000111101101111011011110110","0000111100001111000011110000","0000111110001111100011111000","0000111111111111111111111111","0000101111101011111010111110","0000101011001010110010101100","0000101001111010011110100111","0000101111011011110110111101","0000000010010000100100001001","0000110011001100110011001100","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000011111110111111101111111","0000001111000011110000111100","0000111000101110001011100010","0000011100000111000001110000","0000011100010111000101110001","0000011100100111001001110010","0000101101111011011110110111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111111001111110011111100","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111000111110001111100011","0000101001111010011110100111","0000100111111001111110011111","0000101011111010111110101111","0000111111111111111111111111","0000100010101000101010001010","0000011101000111010001110100","0000101111101011111010111110","0000100011011000110110001101","0000100011111000111110001111","0000110101111101011111010111","0000111110001111100011111000","0000111111011111110111111101","0000111111001111110011111100","0000111110101111101011111010","0000111001001110010011100100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111011111110111111101","0000111100111111001111110011","0000111100001111000011110000","0000110011011100110111001101","0000111111111111111111111111","0000111011101110111011101110","0000111111001111110011111100","0000111010001110100011101000","0000111111111111111111111111","0000111101001111010011110100","0000101100101011001010110010","0000001011100010111000101110","0001000000000000000000000000","0000011100110111001101110011","0000011010010110100101101001","0000010011010100110101001101","0000001110110011101100111011","0000011101000111010001110100","0000111000011110000111100001","0000100110011001100110011001","0000111000111110001111100011","0000111010101110101011101010","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000101100001011000010110000","0000101110111011101110111011","0000111110111111101111111011","0000111101101111011011110110","0000100101111001011110010111","0000011011000110110001101100","0000001000100010001000100010","0000001101100011011000110110","0000011111000111110001111100","0000110000101100001011000010","0000101101111011011110110111","0000110111001101110011011100","0000011011010110110101101101","0000011001100110011001100110","0000011011100110111001101110","0000001001100010011000100110","0001000000000000000000000000","0000000110010001100100011001","0000100010001000100010001000","0000011001100110011001100110","0000101000001010000010100000","0000100101101001011010010110","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111010001110100011101000","0000110110011101100111011001","0000111000111110001111100011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111100111111001111110011","0000111110011111100111111001","0000111110011111100111111001","0000111101111111011111110111","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111111011111110111111101","0000111110101111101011111010","0000111100011111000111110001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000101000011010000110100001","0000111101101111011011110110","0000101010111010101110101011","0000111110011111100111111001","0000110010001100100011001000","0000000110010001100100011001","0000001010110010101100101011","0000100100001001000010010000","0000100100011001000110010001","0000101111011011110110111101","0000101001101010011010100110","0000110111101101111011011110","0000110000011100000111000001","0000011000100110001001100010","0000001011110010111100101111","0000001010000010100000101000","0001000000000000000000000000","0000001111110011111100111111","0000100100011001000110010001","0000101011011010110110101101","0000101110111011101110111011","0000110001111100011111000111","0000110100111101001111010011","0000110101011101010111010101","0000111001011110010111100101","0000101111011011110110111101","0000000100000001000000010000","0000001001100010011000100110","0000000011100000111000001110","0000010000110100001101000011","0000010101000101010001010100","0000011110000111100001111000","0000110101111101011111010111","0000111011011110110111101101","0000111100001111000011110000","0000110110001101100011011000","0000110010101100101011001010","0000100100101001001010010010","0000100111011001110110011101","0000010001010100010101000101","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101011111010111110101","0000111011101110111011101110","0000000101110001011100010111","0000010101000101010001010100","0000010111010101110101011101","0000100001001000010010000100","0000100001011000010110000101","0000111100111111001111110011","0000111100101111001011110010","0000111011111110111111101111","0000111111001111110011111100","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111011101110111011101110","0000110000001100000011000000","0000110000001100000011000000","0000101011101010111010101110","0000111111111111111111111111","0000111000011110000111100001","0000101010001010100010101000","0000101111001011110010111100","0000101101101011011010110110","0000111000011110000111100001","0000110011011100110111001101","0000110110101101101011011010","0000111100101111001011110010","0000111000011110000111100001","0000111111111111111111111111","0000111100101111001011110010","0000111110111111101111111011","0000111101111111011111110111","0000111100001111000011110000","0000111111111111111111111111","0000111100111111001111110011","0000111110011111100111111001","0000111111111111111111111111","0000111010101110101011101010","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000101111111011111110111111","0000100101101001011010010110","0000000000110000001100000011","0000001010110010101100101011","0000010101000101010001010100","0000010010100100101001001010","0000001111000011110000111100","0000001001100010011000100110","0000100100011001000110010001","0000011110000111100001111000","0000110011001100110011001100","0000110011101100111011001110","0000111100011111000111110001","0000100111101001111010011110","0000011111100111111001111110","0000111100111111001111110011","0000111100011111000111110001","0000111111111111111111111111","0000100001101000011010000110","0000100011101000111010001110","0000010001110100011101000111","0000001100010011000100110001","0000110100001101000011010000","0000101011011010110110101101","0000101000101010001010100010","0000101101011011010110110101","0000100111011001110110011101","0000010010110100101101001011","0000010001000100010001000100","0000010111110101111101011111","0000001101000011010000110100","0000001110000011100000111000","0000001111000011110000111100","0000100001001000010010000100","0001000000000000000000000000","0000101011001010110010101100","0000110001101100011011000110","0000111111011111110111111101","0000111101101111011011110110","0000111110101111101011111010","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111001111110011111100","0000111010111110101111101011","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101111111011111110111","0000111111011111110111111101","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111110001111100011111000","0000111010111110101111101011","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111110111111101111111011","0000111111001111110011111100","0000111110111111101111111011","0000111011101110111011101110","0000101101011011010110110101","0000100110011001100110011001","0000111001111110011111100111","0000110001011100010111000101","0000111111111111111111111111","0000101110001011100010111000","0000000111010001110100011101","0001000000000000000000000000","0000100110111001101110011011","0000011111110111111101111111","0000011110110111101101111011","0000101011101010111010101110","0000110101011101010111010101","0000100111001001110010011100","0000011000110110001101100011","0000100000101000001010000010","0000001011110010111100101111","0000010100110101001101010011","0000011000100110001001100010","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000110111011101110111011101","0000010000000100000001000000","0000000111010001110100011101","0000010100010101000101010001","0000010110110101101101011011","0000101011101010111010101110","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000101100011011000110110001","0000111100101111001011110010","0000110010111100101111001011","0000000001000000010000000100","0000101000101010001010100010","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000101101011011010110110101","0001000000000000000000000000","0000011011000110110001101100","0000100000011000000110000001","0000101101011011010110110101","0000111111111111111111111111","0000111011101110111011101110","0000111100101111001011110010","0000111011101110111011101110","0000111010111110101111101011","0000111110001111100011111000","0000111101101111011011110110","0000111110011111100111111001","0000111111111111111111111111","0000111100111111001111110011","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111011111110111111101111","0000111001011110010111100101","0000111101001111010011110100","0000110110011101100111011001","0000110101101101011011010110","0000111111111111111111111111","0000111111111111111111111111","0000110101101101011011010110","0000110110101101101011011010","0000101110001011100010111000","0000110110011101100111011001","0000110101001101010011010100","0000111101001111010011110100","0000111100001111000011110000","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000111101111111011111110111","0000111111111111111111111111","0000111101101111011011110110","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110001111100011111000","0000111101111111011111110111","0000111110111111101111111011","0000111110011111100111111001","0000101101001011010010110100","0000110000001100000011000000","0001000000000000000000000000","0000001001000010010000100100","0000001101100011011000110110","0000010010100100101001001010","0000001010010010100100101001","0000010001000100010001000100","0000010010100100101001001010","0000010011010100110101001101","0000010101010101010101010101","0000100001011000010110000101","0000110011111100111111001111","0000111000111110001111100011","0000111001101110011011100110","0000111111011111110111111101","0000011101010111010101110101","0000100101001001010010010100","0000010101000101010001010100","0001000000000000000000000000","0000110000001100000011000000","0000101000011010000110100001","0000111101001111010011110100","0000011110010111100101111001","0000110100101101001011010010","0000011101110111011101110111","0000011101010111010101110101","0000010001000100010001000100","0000000100110001001100010011","0000000100010001000100010001","0000001110010011100100111001","0000010100110101001101010011","0000010000110100001101000011","0000000010000000100000001000","0000010011010100110101001101","0000111010101110101011101010","0000111111111111111111111111","0000111001111110011111100111","0000111100001111000011110000","0000111111111111111111111111","0000111110101111101011111010","0000111010101110101011101010","0000111111001111110011111100","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111110001111100011111000","0000111111011111110111111101","0000111001011110010111100101","0000111101101111011011110110","0000111111001111110011111100","0000111111001111110011111100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111011001110110011101100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000110010111100101111001011","0000101000101010001010100010","0000100000011000000110000001","0000110101111101011111010111","0000110011101100111011001110","0000111100111111001111110011","0000101001111010011110100111","0000000011010000110100001101","0000010111010101110101011101","0000100101101001011010010110","0000100110101001101010011010","0000011011100110111001101110","0000110001111100011111000111","0000110101111101011111010111","0000110011101100111011001110","0000101111111011111110111111","0000100010111000101110001011","0000001101010011010100110101","0000011001110110011101100111","0000100101101001011010010110","0000110011011100110111001101","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111100111111001111110011","0000111110011111100111111001","0000111101111111011111110111","0000101111001011110010111100","0000010010010100100101001001","0000011101010111010101110101","0000101010101010101010101010","0000100000001000000010000000","0000111111111111111111111111","0000111000101110001011100010","0000100111001001110010011100","0000101111111011111110111111","0000111100001111000011110000","0000101000111010001110100011","0000000100100001001000010010","0000111011101110111011101110","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101101111011011110110","0000111101101111011011110110","0000111100011111000111110001","0000011000000110000001100000","0000000110000001100000011000","0000011101010111010101110101","0000100110001001100010011000","0000111110101111101011111010","0000111111111111111111111111","0000111110011111100111111001","0000110110001101100011011000","0000111101111111011111110111","0000111111111111111111111111","0000110111101101111011011110","0000111001001110010011100100","0000111101011111010111110101","0000111111111111111111111111","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111011011110110111101101","0000111110011111100111111001","0000111100011111000111110001","0000110011001100110011001100","0000110111101101111011011110","0000111111111111111111111111","0000111101011111010111110101","0000111001011110010111100101","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111101001111010011110100","0000111101011111010111110101","0000110100111101001111010011","0000110100111101001111010011","0000100111001001110010011100","0000100110101001101010011010","0000100000011000000110000001","0000011110000111100001111000","0000100000001000000010000000","0000101000111010001110100011","0000101110011011100110111001","0000110110111101101111011011","0000111111111111111111111111","0000111101011111010111110101","0000111001001110010011100100","0000111111111111111111111111","0000111110101111101011111010","0000111111011111110111111101","0000101110001011100010111000","0000110100101101001011010010","0000001010010010100100101001","0000000001110000011100000111","0000100010101000101010001010","0000100000011000000110000001","0000010001100100011001000110","0000001011000010110000101100","0000100000011000000110000001","0000100011011000110110001101","0000010110110101101101011011","0000100110001001100010011000","0000100101111001011110010111","0000100111101001111010011110","0000011010110110101101101011","0000100000101000001010000010","0000010111000101110001011100","0000010111000101110001011100","0000101010101010101010101010","0000101101001011010010110100","0000110111111101111111011111","0000110011001100110011001100","0000101001011010010110100101","0000100111101001111010011110","0000100001101000011010000110","0000100000101000001010000010","0000001000110010001100100011","0000010000100100001001000010","0000000110000001100000011000","0000001011000010110000101100","0000001111110011111100111111","0000001001110010011100100111","0000001011100010111000101110","0001000000000000000000000000","0000111000101110001011100010","0000111111001111110011111100","0000111001001110010011100100","0000111100011111000111110001","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111111111111111111111111","0000111110011111100111111001","0000111100111111001111110011","0000111110001111100011111000","0000111101011111010111110101","0000111010011110100111101001","0000111010001110100011101000","0000111100011111000111110001","0000110010111100101111001011","0000110100001101000011010000","0000110011011100110111001101","0000110101001101010011010100","0000110011001100110011001100","0000110001101100011011000110","0000111000101110001011100010","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111001101110011011100110","0000101111011011110110111101","0000100100011001000110010001","0000100001011000010110000101","0000101100101011001010110010","0000110000101100001011000010","0000110010101100101011001010","0000010000110100001101000011","0000001011000010110000101100","0000101100001011000010110000","0000101110011011100110111001","0000100100001001000010010000","0000100011111000111110001111","0000100001011000010110000101","0000101001101010011010100110","0000110011011100110111001101","0000101111101011111010111110","0000101000111010001110100011","0000011111100111111001111110","0000011101010111010101110101","0000100001011000010110000101","0000101010001010100010101000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111010111110101111101011","0000111000111110001111100011","0000111111111111111111111111","0000111101001111010011110100","0000111111011111110111111101","0000111110001111100011111000","0000101101001011010010110100","0000100110011001100110011001","0000100000001000000010000000","0000011111100111111001111110","0000100110111001101110011011","0000111011101110111011101110","0000110010111100101111001011","0000101001101010011010100110","0000101100011011000110110001","0000110000101100001011000010","0000100001101000011010000110","0000110001101100011011000110","0000111111111111111111111111","0000111101101111011011110110","0000111100011111000111110001","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000110010011100100111001001","0000000011110000111100001111","0000010011110100111101001111","0000100011111000111110001111","0000111100101111001011110010","0000111111111111111111111111","0000111101111111011111110111","0000110110111101101111011011","0000111100101111001011110010","0000111101111111011111110111","0000110111101101111011011110","0000111000101110001011100010","0000111010001110100011101000","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000111111111111111111111111","0000111100001111000011110000","0000111111101111111011111110","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111110111111101111111011","0000110101011101010111010101","0000111101011111010111110101","0000111111111111111111111111","0000111011101110111011101110","0000111100101111001011110010","0000101110111011101110111011","0000101010101010101010101010","0000011011100110111001101110","0000010110000101100001011000","0000100010111000101110001011","0000011010100110101001101010","0000100011101000111010001110","0000100110011001100110011001","0000101011011010110110101101","0000101111101011111010111110","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110001111100011111000","0000111111111111111111111111","0000111100101111001011110010","0000111111011111110111111101","0000111101001111010011110100","0000111010011110100111101001","0000110101001101010011010100","0000111001011110010111100101","0000010001010100010101000101","0000000000110000001100000011","0000101101001011010010110100","0000101011111010111110101111","0000010111010101110101011101","0000010000110100001101000011","0000011000000110000001100000","0000100101011001010110010101","0000100001001000010010000100","0000010111100101111001011110","0000011000000110000001100000","0000010111010101110101011101","0000011000000110000001100000","0000010111000101110001011100","0000011000010110000101100001","0000110110011101100111011001","0000111101101111011011110110","0000101100001011000010110000","0000110101111101011111010111","0000110101101101011011010110","0000100110001001100010011000","0000010100100101001001010010","0000011111000111110001111100","0001000000000000000000000000","0000011001000110010001100100","0000000011000000110000001100","0000001100110011001100110011","0000001101110011011100110111","0000010010100100101001001010","0000001111110011111100111111","0000000100010001000100010001","0000111100011111000111110001","0000111111111111111111111111","0000111001001110010011100100","0000111100111111001111110011","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111100101111001011110010","0000111001101110011011100110","0000110111111101111111011111","0000110111001101110011011100","0000110101011101010111010101","0000110011001100110011001100","0000111000001110000011100000","0000110110111101101111011011","0000110010011100100111001001","0000110011111100111111001111","0000110001111100011111000111","0000101100011011000110110001","0000101101111011011110110111","0000101101001011010010110100","0000111000011110000111100001","0000111101011111010111110101","0000110100001101000011010000","0000100110111001101110011011","0000100000111000001110000011","0000010110110101101101011011","0000010001110100011101000111","0000011001110110011101100111","0000011000000110000001100000","0000011010110110101101101011","0001000000000000000000000000","0000010001110100011101000111","0000110111011101110111011101","0000101101101011011010110110","0000101000111010001110100011","0000100010111000101110001011","0000011110100111101001111010","0000011011010110110101101101","0000100000011000000110000001","0000011110110111101101111011","0000101111101011111010111110","0000110010001100100011001000","0000101011001010110010101100","0000011000000110000001100000","0000100110011001100110011001","0000110000101100001011000010","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111110001111100011111000","0000111111101111111011111110","0000110010111100101111001011","0000101101011011010110110101","0000100000101000001010000010","0000100111001001110010011100","0000011101110111011101110111","0000110110001101100011011000","0000101111001011110010111100","0000101100101011001010110010","0000110011011100110111001101","0000011110110111101101111011","0000011011100110111001101110","0000111101101111011011110110","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000110010111100101111001011","0000001101010011010100110101","0001000000000000000000000000","0000101000001010000010100000","0000111001111110011111100111","0000111111001111110011111100","0000111111001111110011111100","0000111101011111010111110101","0000110100011101000111010001","0000110000011100000111000001","0000111011011110110111101101","0000111111111111111111111111","0000111101111111011111110111","0000110011011100110111001101","0000111101111111011111110111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111011101110111011101110","0000111110011111100111111001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111100011111000111110001","0000101110101011101010111010","0000111000111110001111100011","0000111111111111111111111111","0000110011001100110011001100","0000100011011000110110001101","0000010010000100100001001000","0001000000000000000000000000","0001000000000000000000000000","0000010011010100110101001101","0000101001101010011010100110","0000101101101011011010110110","0000110000001100000011000000","0000110100111101001111010011","0000111000101110001011100010","0000110010101100101011001010","0000110001001100010011000100","0000111000111110001111100011","0000111100001111000011110000","0000111101011111010111110101","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000110100111101001111010011","0000110011001100110011001100","0000011011110110111101101111","0000000001100000011000000110","0000100011101000111010001110","0000101111111011111110111111","0000101101001011010010110100","0000010111000101110001011100","0000010100110101001101010011","0000000100110001001100010011","0000011100010111000101110001","0000010011010100110101001101","0000010110000101100001011000","0000001111000011110000111100","0000101000111010001110100011","0000110001111100011111000111","0000111101101111011011110110","0000110011101100111011001110","0000111111111111111111111111","0000110100011101000111010001","0000110101101101011011010110","0000011110010111100101111001","0000001111010011110100111101","0000010000110100001101000011","0000000000100000001000000010","0000010001000100010001000100","0000000010110000101100001011","0000010001110100011101000111","0000001011110010111100101111","0000010000000100000001000000","0000010101110101011101010111","0000000110000001100000011000","0000111000111110001111100011","0000111111111111111111111111","0000110000001100000011000000","0000110111011101110111011101","0000111100001111000011110000","0000111111111111111111111111","0000111101101111011011110110","0000111011001110110011101100","0000111100111111001111110011","0000111101011111010111110101","0000111010101110101011101010","0000110110001101100011011000","0000110001111100011111000111","0000101110111011101110111011","0000101101011011010110110101","0000110010101100101011001010","0000101110011011100110111001","0000100011001000110010001100","0000100010101000101010001010","0000100111101001111010011110","0000101010101010101010101010","0000101011101010111010101110","0000100011011000110110001101","0000010000110100001101000011","0000010011010100110101001101","0000000101110001011100010111","0001000000000000000000000000","0000000100100001001000010010","0000000011000000110000001100","0001000000000000000000000000","0000001000110010001100100011","0000010110110101101101011011","0000110001111100011111000111","0000101111101011111010111110","0000100001101000011010000110","0000011000000110000001100000","0000011001110110011101100111","0000011110000111100001111000","0000011010110110101101101011","0000011000100110001001100010","0000101100111011001110110011","0000100110111001101110011011","0000010111110101111101011111","0000100010101000101010001010","0000110110001101100011011000","0000011111100111111001111110","0000011110010111100101111001","0000100110111001101110011011","0000111101101111011011110110","0000111110101111101011111010","0000111010101110101011101010","0000111111001111110011111100","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010001110100011101000","0000111011001110110011101100","0000111110011111100111111001","0000110101001101010011010100","0000110101101101011011010110","0000100111001001110010011100","0000100101011001010110010101","0000011111000111110001111100","0000101010001010100010101000","0000100111011001110110011101","0000101110011011100110111001","0000101100011011000110110001","0000010111100101111001011110","0000110001111100011111000111","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000111010101110101011101010","0000111010011110100111101001","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000100010111000101110001011","0000001001100010011000100110","0000001000010010000100100001","0000100010111000101110001011","0000111111011111110111111101","0000111111101111111011111110","0000111001111110011111100111","0000111111111111111111111111","0000111011001110110011101100","0000100110001001100010011000","0000110010011100100111001001","0000111111111111111111111111","0000110110011101100111011001","0000101100111011001110110011","0000111101111111011111110111","0000111010101110101011101010","0000111000111110001111100011","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110111111101111111011","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111011101110111011101110","0000100101101001011010010110","0000110010011100100111001001","0000101010011010100110101001","0000100000101000001010000010","0000000101000001010000010100","0000000010000000100000001000","0000001100100011001000110010","0000011110100111101001111010","0000100000101000001010000010","0000101010111010101110101011","0000110011001100110011001100","0000110000001100000011000000","0000110000101100001011000010","0000110100111101001111010011","0000110100011101000111010001","0000110110101101101011011010","0000110111101101111011011110","0000111100101111001011110010","0000111111101111111011111110","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111001111110011111100","0000111110101111101011111010","0000111100011111000111110001","0000111101011111010111110101","0000111111111111111111111111","0000101111101011111010111110","0000111100111111001111110011","0000101100001011000010110000","0000000001100000011000000110","0000001110010011100100111001","0000101111111011111110111111","0000111000001110000011100000","0000100011111000111110001111","0000101000011010000110100001","0000010110100101101001011010","0000011111110111111101111111","0000101010001010100010101000","0000011111010111110101111101","0000110100011101000111010001","0000110101001101010011010100","0000111011011110110111101101","0000111010101110101011101010","0000111111111111111111111111","0000111100001111000011110000","0000110111111101111111011111","0000011011010110110101101101","0000010000000100000001000000","0001000000000000000000000000","0000000100100001001000010010","0000010110000101100001011000","0000000011000000110000001100","0000010110100101101001011010","0000011000010110000101100001","0000010001000100010001000100","0000001011000010110000101100","0000010100010101000101010001","0000101000011010000110100001","0000101110101011101010111010","0000100111001001110010011100","0000111000101110001011100010","0000111011111110111111101111","0000111111111111111111111111","0000111011101110111011101110","0000111000001110000011100000","0000111011001110110011101100","0000101111111011111110111111","0000101111101011111010111110","0000100000101000001010000010","0000100011011000110110001101","0000101000111010001110100011","0000101011101010111010101110","0000110100101101001011010010","0000110111111101111111011111","0000111001111110011111100111","0000111011111110111111101111","0000110100101101001011010010","0000011011110110111101101111","0000000101000001010000010100","0001000000000000000000000000","0001000000000000000000000000","0000000111110001111100011111","0000010110110101101101011011","0000010010100100101001001010","0000011000110110001101100011","0000101110011011100110111001","0000110110101101101011011010","0000111111111111111111111111","0000111111111111111111111111","0000110101001101010011010100","0000101111111011111110111111","0000101110001011100010111000","0000100011001000110010001100","0000010110110101101101011011","0000010100010101000101010001","0000010111010101110101011101","0000011001000110010001100100","0000010110100101101001011010","0000011011010110110101101101","0000100110111001101110011011","0000100110001001100010011000","0000100100011001000110010001","0000111000001110000011100000","0000100100111001001110010011","0000101100011011000110110001","0000111101001111010011110100","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111100101111001011110010","0000110100011101000111010001","0000111110011111100111111001","0000111111101111111011111110","0000110001111100011111000111","0000101111101011111010111110","0000101001001010010010100100","0000010101110101011101010111","0000100101101001011010010110","0000011100010111000101110001","0000101001111010011110100111","0000011111100111111001111110","0000101011001010110010101100","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111110001111100011111000","0000111101001111010011110100","0000110010101100101011001010","0000011110010111100101111001","0000001101100011011000110110","0000010110110101101101011011","0000100011001000110010001100","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111000101110001011100010","0000001001110010011100100111","0000100010011000100110001001","0000101110111011101110111011","0000110001001100010011000100","0000101111111011111110111111","0000111101001111010011110100","0000111111111111111111111111","0000110011111100111111001111","0000111111111111111111111111","0000111111001111110011111100","0000111010111110101111101011","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111110101111101011111010","0000100110111001101110011011","0000110011111100111111001111","0000100001101000011010000110","0000011010110110101101101011","0001000000000000000000000000","0000001101000011010000110100","0000011110010111100101111001","0000100001011000010110000101","0000011111100111111001111110","0000101010111010101110101011","0000110100011101000111010001","0000111000101110001011100010","0000110010111100101111001011","0000110011101100111011001110","0000111010101110101011101010","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111100111111001111110011","0000111101011111010111110101","0000111111001111110011111100","0000111111111111111111111111","0000111000101110001011100010","0000111001111110011111100111","0000111110111111101111111011","0000101101111011011110110111","0000100000101000001010000010","0000011001000110010001100100","0000100100011001000110010001","0000101011101010111010101110","0000100101001001010010010100","0000101101101011011010110110","0000100110001001100010011000","0000101110111011101110111011","0000011110110111101101111011","0000101111101011111010111110","0000111100101111001011110010","0000100110001001100010011000","0000111110101111101011111010","0000111001011110010111100101","0000111111111111111111111111","0000110011101100111011001110","0000011000010110000101100001","0000001100100011001000110010","0000001100100011001000110010","0000001010110010101100101011","0000011101010111010101110101","0000000001110000011100000111","0000010100100101001001010010","0000010010000100100001001000","0000001110100011101000111010","0000011100110111001101110011","0000001111110011111100111111","0000010111100101111001011110","0000011011110110111101101111","0000011111010111110101111101","0000111100101111001011110010","0000111111111111111111111111","0000111101111111011111110111","0000101111011011110110111101","0000110111101101111011011110","0000100010011000100110001001","0000110011011100110111001101","0000001111110011111100111111","0000011000010110000101100001","0000100101011001010110010101","0000101010111010101110101011","0000101111111011111110111111","0000101111111011111110111111","0000100110111001101110011011","0000011100100111001001110010","0000001101000011010000110100","0001000000000000000000000000","0000000101010001010100010101","0000010110110101101101011011","0000100000011000000110000001","0000100111011001110110011101","0000100101111001011110010111","0000101011111010111110101111","0000110011111100111111001111","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000110111011101110111011101","0000110101111101011111010111","0000110110011101100111011001","0000110101111101011111010111","0000110101011101010111010101","0000110010001100100011001000","0000101011011010110110101101","0000100100001001000010010000","0000100000001000000010000000","0000010011010100110101001101","0000001011110010111100101111","0000101100101011001010110010","0000101101111011011110110111","0000101001111010011110100111","0000011011010110110101101101","0000110101001101010011010100","0000111110001111100011111000","0000111110011111100111111001","0000111111001111110011111100","0000111110011111100111111001","0000111010101110101011101010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000110110011101100111011001","0000110110101101101011011010","0000111010001110100011101000","0000111010111110101111101011","0000110111101101111011011110","0000100000001000000010000000","0000101000001010000010100000","0000100100101001001010010010","0000100101011001010110010101","0000100000001000000010000000","0000010101000101010001010100","0000011000000110000001100000","0000111011111110111111101111","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111111101111111011111110","0000110100111101001111010011","0000011101100111011001110110","0000000010010000100100001001","0000010111100101111001011110","0000101011001010110010101100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000110101101101011011010110","0000010100110101001101010011","0000100011011000110110001101","0000101011011010110110101101","0000101111011011110110111101","0000110010111100101111001011","0000110111101101111011011110","0000111101101111011011110110","0000101110001011100010111000","0000110101001101010011010100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101101101011011010110110","0000100001111000011110000111","0000010111100101111001011110","0000011101010111010101110101","0000000100000001000000010000","0000010001010100010101000101","0000100010101000101010001010","0000100011001000110010001100","0000100000011000000110000001","0000100010111000101110001011","0000101000001010000010100000","0000110010101100101011001010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000110101111101011111010111","0000111010011110100111101001","0000111010001110100011101000","0000110110111101101111011011","0000111101111111011111110111","0000111001001110010011100100","0000110010101100101011001010","0000101001011010010110100101","0000011100100111001001110010","0000011011000110110001101100","0000100010001000100010001000","0000110010111100101111001011","0000011010110110101101101011","0000011110000111100001111000","0000101100011011000110110001","0000110010011100100111001001","0000101110101011101010111010","0000111001011110010111100101","0000111100001111000011110000","0000111110101111101011111010","0000101111001011110010111100","0000101111101011111010111110","0000001111000011110000111100","0000001010010010100100101001","0000001000110010001100100011","0000010001000100010001000100","0000010100000101000001010000","0001000000000000000000000000","0000001011110010111100101111","0000000110000001100000011000","0000001101000011010000110100","0000011111110111111101111111","0000001010010010100100101001","0000001110110011101100111011","0000010101100101011001010110","0000011010100110101001101010","0000110111011101110111011101","0000111011001110110011101100","0000100111011001110110011101","0000001110110011101100111011","0000010110100101101001011010","0000110101111101011111010111","0000011000000110000001100000","0000011001110110011101100111","0000011100010111000101110001","0000101011101010111010101110","0000101000101010001010100010","0000011000010110000101100001","0000000001010000010100000101","0000000011100000111000001110","0000001111010011110100111101","0000011111000111110001111100","0000101110111011101110111011","0000111111001111110011111100","0000111111111111111111111111","0000111010001110100011101000","0000111010111110101111101011","0000111100111111001111110011","0000111100011111000111110001","0000111110111111101111111011","0000111110001111100011111000","0000111011001110110011101100","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000110100111101001111010011","0000101011001010110010101100","0000100001011000010110000101","0000100100111001001110010011","0000101001001010010010100100","0000100101101001011010010110","0000100111111001111110011111","0000001010100010101000101010","0000000110110001101100011011","0000100111001001110010011100","0000011010010110100101101001","0000111011001110110011101100","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110110101101101011011010","0000111101101111011011110110","0000110111101101111011011110","0000111111111111111111111111","0000111110101111101011111010","0000010101100101011001010110","0000011001110110011101100111","0000100000011000000110000001","0000100100011001000110010001","0000100001011000010110000101","0000000001010000010100000101","0000101010111010101110101011","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111001111110011111100","0000110011011100110111001101","0000100101011001010110010101","0000000010100000101000001010","0000011010110110101101101011","0000101111101011111010111110","0000111100001111000011110000","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111110001111100011111000","0000010111110101111101011111","0000011111000111110001111100","0000101000111010001110100011","0000101001001010010010100100","0000101001001010010010100100","0000101100001011000010110000","0000101000101010001010100010","0000100101011001010110010101","0000100011111000111110001111","0000101110111011101110111011","0000110001111100011111000111","0000011111010111110101111101","0000100000101000001010000010","0000011001110110011101100111","0000100111111001111110011111","0000001010000010100000101000","0000011100100111001001110010","0000101001011010010110100101","0000100011011000110110001101","0000010011010100110101001101","0000100101111001011110010111","0000110001011100010111000101","0000101101101011011010110110","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111100111111001111110011","0000111110001111100011111000","0000111011001110110011101100","0000111111111111111111111111","0000111001011110010111100101","0000110110101101101011011010","0000111011101110111011101110","0000111111111111111111111111","0000111111011111110111111101","0000111101101111011011110110","0000111101111111011111110111","0000110110111101101111011011","0000101111011011110110111101","0000101010111010101110101011","0000110000001100000011000000","0000110100111101001111010011","0000110011001100110011001100","0000101110101011101010111010","0000101001101010011010100110","0000101000101010001010100010","0000010111100101111001011110","0000001111110011111100111111","0000010000010100000101000001","0000011010000110100001101000","0000011111100111111001111110","0000101010111010101110101011","0000101000111010001110100011","0000101110001011100010111000","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111010101110101011101010","0000011101000111010001110100","0000001110100011101000111010","0000011101000111010001110100","0000000110000001100000011000","0000001000000010000000100000","0000001001000010010000100100","0000000101010001010100010101","0000001000010010000100100001","0000001010110010101100101011","0000000101000001010000010100","0000011010010110100101101001","0000010100000101000001010000","0000000110110001101100011011","0000001010000010100000101000","0000010011000100110001001100","0000100000111000001110000011","0000010111000101110001011100","0000001110100011101000111010","0000010100010101000101010001","0000101011111010111110101111","0000100110011001100110011001","0000011001110110011101100111","0000011001110110011101100111","0000100110111001101110011011","0000010011110100111101001111","0000001110110011101100111011","0000100011111000111110001111","0000011100110111001101110011","0000101100001011000010110000","0000110111011101110111011101","0000111101001111010011110100","0000111111111111111111111111","0000111111001111110011111100","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101101111011011110110","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111010011110100111101001","0000110100101101001011010010","0000101000011010000110100001","0000011011100110111001101110","0000011011110110111101101111","0000100001101000011010000110","0000100011111000111110001111","0000001111010011110100111101","0000001000100010001000100010","0000011011100110111001101110","0000110111011101110111011101","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111011101110111011101110","0000111101001111010011110100","0000110011001100110011001100","0000111000011110000111100001","0000110010011100100111001001","0000111111111111111111111111","0000110010101100101011001010","0000011000100110001001100010","0000110101111101011111010111","0000100111001001110010011100","0000011111000111110001111100","0000000001000000010000000100","0000011111100111111001111110","0000111111101111111011111110","0000111111111111111111111111","0000111001101110011011100110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000101100101011001010110010","0000100011101000111010001110","0001000000000000000000000000","0000010111110101111101011111","0000110000101100001011000010","0000111101001111010011110100","0000111110001111100011111000","0000111111001111110011111100","0000111111001111110011111100","0000111010001110100011101000","0000100010001000100010001000","0001000000000000000000000000","0000001011000010110000101100","0000011100110111001101110011","0000011100010111000101110001","0000100000111000001110000011","0000101001111010011110100111","0000101000101010001010100010","0000011000010110000101100001","0000010011000100110001001100","0000011000010110000101100001","0000010001100100011001000110","0000101011001010110010101100","0000011001100110011001100110","0000001111000011110000111100","0000100011111000111110001111","0000101111111011111110111111","0000011011110110111101101111","0000011100000111000001110000","0000110000111100001111000011","0000110010011100100111001001","0000110101011101010111010101","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111010001110100011101000","0000111000001110000011100000","0000110000111100001111000011","0000100111011001110110011101","0000100110101001101010011010","0000100110011001100110011001","0000100110101001101010011010","0000100111011001110110011101","0000101011111010111110101111","0000110101011101010111010101","0000111110001111100011111000","0000111011001110110011101100","0000101011011010110110101101","0000100010001000100010001000","0000100100001001000010010000","0000100111101001111010011110","0000110111001101110011011100","0000100100001001000010010000","0000011001110110011101100111","0000100001011000010110000101","0000101001111010011110100111","0000100011101000111010001110","0000100001111000011110000111","0000011110000111100001111000","0000011111100111111001111110","0000100010111000101110001011","0000100001001000010010000100","0000101001001010010010100100","0000110100101101001011010010","0000110011111100111111001111","0000111000111110001111100011","0000101000011010000110100001","0000011111110111111101111111","0000010000010100000101000001","0000011110110111101101111011","0001000000000000000000000000","0000011011110110111101101111","0000001001110010011100100111","0000000100110001001100010011","0000000110100001101000011010","0000011001010110010101100101","0000011110110111101101111011","0000000001000000010000000100","0000010001110100011101000111","0000000110110001101100011011","0000001000010010000100100001","0000001000010010000100100001","0000001000010010000100100001","0000000010000000100000001000","0000001010000010100000101000","0000011111110111111101111111","0000011000000110000001100000","0000010100100101001001010010","0000010100100101001001010010","0000011000010110000101100001","0000011101010111010101110101","0000100000111000001110000011","0000100111101001111010011110","0000101001111010011110100111","0000110110001101100011011000","0000111101101111011011110110","0000111110111111101111111011","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111100011111000111110001","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111011001110110011101100","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111011011110110111101101","0000111100111111001111110011","0000111111111111111111111111","0000111101101111011011110110","0000101111101011111010111110","0000111111111111111111111111","0000111001001110010011100100","0000100101111001011110010111","0000100001001000010010000100","0000011010010110100101101001","0000100111001001110010011100","0001000000000000000000000000","0000010001110100011101000111","0000110011011100110111001101","0000111101011111010111110101","0000111101001111010011110100","0000111101011111010111110101","0000111111001111110011111100","0000111110011111100111111001","0000111111101111111011111110","0000111101011111010111110101","0000110111011101110111011101","0000110111111101111111011111","0000011100100111001001110010","0000101001011010010110100101","0000101100101011001010110010","0000110001001100010011000100","0000100000101000001010000010","0000101101001011010010110100","0000101010101010101010101010","0000100101001001010010010100","0001000000000000000000000000","0000011111100111111001111110","0000111111111111111111111111","0000111111011111110111111101","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110011111100111111001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111101011111010111110101","0000101111011011110110111101","0000100101011001010110010101","0000000010110000101100001011","0000011100000111000001110000","0000100110101001101010011010","0000111010011110100111101001","0000111011111110111111101111","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000101100101011001010110010","0000010010100100101001001010","0000000101000001010000010100","0000010100000101000001010000","0000011010100110101001101010","0000011000110110001101100011","0000010111000101110001011100","0000100000111000001110000011","0000011001010110010101100101","0000010111000101110001011100","0000011010010110100101101001","0000111111011111110111111101","0000000101100001011000010110","0000011100110111001101110011","0000110101101101011011010110","0000011111010111110101111101","0000010011010100110101001101","0000110000011100000111000001","0000011111110111111101111111","0000101101101011011010110110","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111010101110101011101010","0000110101001101010011010100","0000110101001101010011010100","0000111100011111000111110001","0000111010101110101011101010","0000101100111011001110110011","0000100111001001110010011100","0000100000011000000110000001","0000011010110110101101101011","0000010101100101011001010110","0000010000110100001101000011","0000001111100011111000111110","0000010000100100001001000010","0000011100010111000101110001","0000010101100101011001010110","0000011100010111000101110001","0000011011110110111101101111","0000011100100111001001110010","0000110111101101111011011110","0000011101100111011001110110","0000011011000110110001101100","0000011101000111010001110100","0000100101101001011010010110","0000011101010111010101110101","0000101100111011001110110011","0000100000101000001010000010","0000011100010111000101110001","0000100100101001001010010010","0000100000101000001010000010","0000011100110111001101110011","0000100000001000000010000000","0000101010011010100110101001","0000100011011000110110001101","0000010100010101000101010001","0000011000010110000101100001","0000011111000111110001111100","0000000001010000010100000101","0000001010000010100000101000","0000010100000101000001010000","0000001010000010100000101000","0000000100010001000100010001","0000001010110010101100101011","0000010111110101111101011111","0000011001100110011001100110","0001000000000000000000000000","0000000001010000010100000101","0000000111010001110100011101","0000001100100011001000110010","0000001000010010000100100001","0000001001010010010100100101","0000010000000100000001000000","0000010110110101101101011011","0000011011100110111001101110","0000010110110101101101011011","0000011100000111000001110000","0000100000001000000010000000","0000100010011000100110001001","0000100011011000110110001101","0000101011001010110010101100","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110010011100100111001001","0000101001011010010110100101","0000111110101111101011111010","0000111011101110111011101110","0000011110110111101101111011","0000010111110101111101011111","0000101001001010010010100100","0000000110000001100000011000","0000000011100000111000001110","0000110001111100011111000111","0000111011011110110111101101","0000111100101111001011110010","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111111011111110111111101","0000101111001011110010111100","0000101100011011000110110001","0000010111100101111001011110","0000100000001000000010000000","0000011000010110000101100001","0000110011001100110011001100","0000111111101111111011111110","0000101101111011011110110111","0000101010111010101110101011","0000000100010001000100010001","0000011010000110100001101000","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111011111110111111101","0000111011101110111011101110","0000100110011001100110011001","0000011111100111111001111110","0000000101000001010000010100","0000100001011000010110000101","0000100001111000011110000111","0000101011111010111110101111","0000111000011110000111100001","0000111010101110101011101010","0000111110011111100111111001","0000111111111111111111111111","0000111110101111101011111010","0000100110111001101110011011","0000000010100000101000001010","0000000000100000001000000010","0000100000111000001110000011","0000101000101010001010100010","0000100000011000000110000001","0000100011011000110110001101","0000100111101001111010011110","0000101000001010000010100000","0000010110000101100001011000","0000000011100000111000001110","0000100010001000100010001000","0000100110101001101010011010","0000010110000101100001011000","0000001110010011100100111001","0000010010010100100101001001","0000101011001010110010101100","0000111001001110010011100100","0000111111101111111011111110","0000111111111111111111111111","0000111110011111100111111001","0000111001111110011111100111","0000111100011111000111110001","0000111101001111010011110100","0000111110011111100111111001","0000111111011111110111111101","0000110100111101001111010011","0000110101001101010011010100","0000011100000111000001110000","0000001001100010011000100110","0000001011110010111100101111","0000010000110100001101000011","0000001101010011010100110101","0000001001100010011000100110","0000001011010010110100101101","0000001111100011111000111110","0000000110100001101000011010","0001000000000000000000000000","0001000000000000000000000000","0000000010110000101100001011","0000011001000110010001100100","0000010000110100001101000011","0000010111000101110001011100","0000100000011000000110000001","0000100101101001011010010110","0000001111100011111000111110","0000011001010110010101100101","0000011001000110010001100100","0000010011110100111101001111","0000001111010011110100111101","0000011000000110000001100000","0000100001001000010010000100","0000011001000110010001100100","0000011111100111111001111110","0000100001101000011010000110","0000100111001001110010011100","0000010110110101101101011011","0000011001010110010101100101","0001000000000000000000000000","0000001001100010011000100110","0000010100010101000101010001","0000000101110001011100010111","0000000011110000111100001111","0000001001010010010100100101","0000001100000011000000110000","0000010101100101011001010110","0000000100100001001000010010","0000001010010010100100101001","0000000001000000010000000100","0000000000110000001100000011","0000010010000100100001001000","0000011110010111100101111001","0000100000001000000010000000","0000100010101000101010001010","0000100101001001010010010100","0000011101010111010101110101","0000100001111000011110000111","0000011100010111000101110001","0000101000011010000110100001","0000111000111110001111100011","0000111111111111111111111111","0000111011111110111111101111","0000111100001111000011110000","0000111111111111111111111111","0000111100101111001011110010","0000111110101111101011111010","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111111001111110011111100","0000111000001110000011100000","0000110001111100011111000111","0000110000011100000111000001","0000101010001010100010101000","0000101001111010011110100111","0000101111101011111010111110","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111101111111011111110111","0000111110011111100111111001","0000100111011001110110011101","0000101101011011010110110101","0000111111111111111111111111","0000101010001010100010101000","0000010000110100001101000011","0000100010011000100110001001","0001000000000000000000000000","0000011011010110110101101101","0000100100101001001010010010","0000110101101101011011010110","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111011011110110111101101","0000100011111000111110001111","0000100110101001101010011010","0000010010100100101001001010","0000011000110110001101100011","0000110010011100100111001001","0000110111001101110011011100","0000110000111100001111000011","0000101010111010101110101011","0001000000000000000000000000","0000100010001000100010001000","0000111001011110010111100101","0000111111011111110111111101","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111110011111100111111001","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000100111001001110010011100","0000010011010100110101001101","0001000000000000000000000000","0000010011110100111101001111","0000100110111001101110011011","0000100000101000001010000010","0000101111111011111110111111","0000110010111100101111001011","0000110101011101010111010101","0000101100011011000110110001","0000110100111101001111010011","0000101111101011111010111110","0000001110000011100000111000","0001000000000000000000000000","0000000010100000101000001010","0000010001110100011101000111","0000001110000011100000111000","0000011100010111000101110001","0000010111110101111101011111","0000010101110101011101010111","0000001111000011110000111100","0000011001000110010001100100","0000001011110010111100101111","0000001001000010010000100100","0000001001100010011000100110","0000011011000110110001101100","0000110111001101110011011100","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101101111011011110110","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111111101111111011111110","0000110101111101011111010111","0000001111100011111000111110","0000100000001000000010000000","0000101000101010001010100010","0000100100011001000110010001","0000100110101001101010011010","0000110001011100010111000101","0000110010101100101011001010","0000101001101010011010100110","0000100010101000101010001010","0000100100011001000110010001","0000010011000100110001001100","0000011001000110010001100100","0000011000010110000101100001","0000010001100100011001000110","0000001011010010110100101101","0000000001100000011000000110","0000000010000000100000001000","0000001100000011000000110000","0000010000010100000101000001","0000100110101001101010011010","0000011111010111110101111101","0000110110101101101011011010","0000100001011000010110000101","0000011100000111000001110000","0000100100011001000110010001","0000010101010101010101010101","0000010101000101010001010100","0000011111000111110001111100","0000111110101111101011111010","0000101001101010011010100110","0000000001110000011100000111","0000001111100011111000111110","0000001011100010111000101110","0000010001010100010101000101","0000001000110010001100100011","0000001010010010100100101001","0000001010000010100000101000","0000001100000011000000110000","0000001100110011001100110011","0000010101010101010101010101","0000011111000111110001111100","0000001000110010001100100011","0001000000000000000000000000","0000011000100110001001100010","0000101010101010101010101010","0000101000001010000010100000","0000100100101001001010010010","0000100010001000100010001000","0000101001111010011110100111","0000110000011100000111000001","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111111111111111111111","0000111110011111100111111001","0000111111011111110111111101","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000110000111100001111000011","0000101011011010110110101101","0000110010111100101111001011","0000100101001001010010010100","0000100011011000110110001101","0000011010000110100001101000","0000011111000111110001111100","0000011100100111001001110010","0000011000000110000001100000","0000101011111010111110101111","0000111000111110001111100011","0000111111111111111111111111","0000111101101111011011110110","0000111101111111011111110111","0000111101111111011111110111","0000111100111111001111110011","0000111110101111101011111010","0000111101111111011111110111","0000111000101110001011100010","0000100110011001100110011001","0000101011011010110110101101","0000111101001111010011110100","0000101000111010001110100011","0000010100100101001001010010","0000010010110100101101001011","0000000110000001100000011000","0000100001111000011110000111","0000010000010100000101000001","0000101100011011000110110001","0000111010101110101011101010","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000110001011100010111000101","0000010110100101101001011010","0000011101010111010101110101","0000100010011000100110001001","0000010011110100111101001111","0000110010001100100011001000","0000111110101111101011111010","0000100101111001011110010111","0001000000000000000000000000","0000100100101001001010010010","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111011011110110111101101","0000111100111111001111110011","0000111111111111111111111111","0000110111001101110011011100","0000011110110111101101111011","0000000111110001111100011111","0001000000000000000000000000","0000010100110101001101010011","0000011011100110111001101110","0000100100011001000110010001","0000101101001011010010110100","0000101101101011011010110110","0000100100111001001110010011","0000100101101001011010010110","0000011011010110110101101101","0000001011100010111000101110","0000010100010101000101010001","0000000110000001100000011000","0000000001000000010000000100","0000000111010001110100011101","0001000000000000000000000000","0000000110010001100100011001","0001000000000000000000000000","0000100001111000011110000111","0000101111111011111110111111","0000011101100111011001110110","0000010000100100001001000010","0000011100100111001001110010","0000111111001111110011111100","0000111011111110111111101111","0000111101011111010111110101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111110011111100111111001","0000110011101100111011001110","0000100111001001110010011100","0000100110111001101110011011","0000100000011000000110000001","0000100100011001000110010001","0000110010001100100011001000","0000110110111101101111011011","0000110001111100011111000111","0000110011101100111011001110","0000111100111111001111110011","0000111001101110011011100110","0000110100111101001111010011","0000111000101110001011100010","0000011110010111100101111001","0000110001111100011111000111","0000101010111010101110101011","0000111001011110010111100101","0000110001011100010111000101","0000011111000111110001111100","0000011000110110001101100011","0001000000000000000000000000","0000000000110000001100000011","0000000011100000111000001110","0000010111000101110001011100","0000011100110111001101110011","0000011111010111110101111101","0000011001110110011101100111","0000101111001011110010111100","0000101100101011001010110010","0000101010111010101110101011","0000010100010101000101010001","0000010000100100001001000010","0000011001100110011001100110","0000011111110111111101111111","0000010101010101010101010101","0000011001100110011001100110","0001000000000000000000000000","0000001000100010001000100010","0000001100100011001000110010","0000011100110111001101110011","0000010110000101100001011000","0000101000111010001110100011","0000011000010110000101100001","0000010100110101001101010011","0000011011100110111001101110","0000011011100110111001101110","0000010001110100011101000111","0000000011100000111000001110","0001000000000000000000000000","0000010010100100101001001010","0000011101100111011001110110","0000100110111001101110011011","0000110010001100100011001000","0000111100011111000111110001","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111011111110111111101","0000110011101100111011001110","0000101010101010101010101010","0000110101001101010011010100","0000110111111101111111011111","0000100110111001101110011011","0000110000111100001111000011","0000100110111001101110011011","0000001111110011111100111111","0001000000000000000000000000","0000010011100100111001001110","0000011001010110010101100101","0000011101000111010001110100","0000001000110010001100100011","0000100110111001101110011011","0000111111111111111111111111","0000111111011111110111111101","0000111101001111010011110100","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000101011011010110110101101","0000101110011011100110111001","0000110101111101011111010111","0000100111011001110110011101","0000011110010111100101111001","0000011101100111011001110110","0000000000100000001000000010","0000010011010100110101001101","0000100011011000110110001101","0000011101110111011101110111","0000010111010101110101011101","0000101100001011000010110000","0000111111111111111111111111","0000111111001111110011111100","0000110100111101001111010011","0000101011111010111110101111","0000011100100111001001110010","0000011011110110111101101111","0000011000110110001101100011","0000010011110100111101001111","0000100011101000111010001110","0000110110001101100011011000","0000001111110011111100111111","0000000100110001001100010011","0000110100111101001111010011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000110111101101111011011110","0000100101001001010010010100","0000000001000000010000000100","0000000000010000000100000001","0000000111110001111100011111","0000100010101000101010001010","0000110101011101010111010101","0000110111101101111011011110","0000010110110101101101011011","0000001010000010100000101000","0000101101011011010110110101","0000101011111010111110101111","0000100101001001010010010100","0000001111100011111000111110","0000010101000101010001010100","0000001100110011001100110011","0000011001010110010101100101","0000001100100011001000110010","0000010011010100110101001101","0000011111110111111101111111","0000100001111000011110000111","0000000101000001010000010100","0000001101110011011100110111","0000100110111001101110011011","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000110010011100100111001001","0000101110111011101110111011","0000101111001011110010111100","0000100110101001101010011010","0000100101101001011010010110","0000100110001001100010011000","0000101011101010111010101110","0000110110111101101111011011","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111100101111001011110010","0000111010111110101111101011","0000111101011111010111110101","0000100110101001101010011010","0000110011101100111011001110","0000110101001101010011010100","0000110101101101011011010110","0000101110101011101010111010","0000111000011110000111100001","0000101000001010000010100000","0000011110110111101101111011","0000010101110101011101010111","0000010011110100111101001111","0000001000100010001000100010","0000000011010000110100001101","0001000000000000000000000000","0000000100100001001000010010","0000001101100011011000110110","0000011010110110101101101011","0000100100011001000110010001","0000100011011000110110001101","0000101001001010010010100100","0000100100111001001110010011","0000010010010100100101001001","0000010001010100010101000101","0000011000000110000001100000","0000001100100011001000110010","0000010100000101000001010000","0000100101101001011010010110","0000001011010010110100101101","0000100010001000100010001000","0000001110110011101100111011","0000100000001000000010000000","0000100100001001000010010000","0000011100110111001101110011","0000100000111000001110000011","0000101101111011011110110111","0000110011111100111111001111","0000110001101100011011000110","0000101111101011111010111110","0000110100001101000011010000","0000111010011110100111101001","0000110111101101111011011110","0000111011111110111111101111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001111110011111100111","0000110110001101100011011000","0000111101101111011011110110","0000111100101111001011110010","0000111001111110011111100111","0000111111111111111111111111","0000100101011001010110010101","0000000001100000011000000110","0000011101010111010101110101","0000111001011110010111100101","0000111111111111111111111111","0000111100011111000111110001","0000110101101101011011010110","0000110101001101010011010100","0000101111111011111110111111","0000101011001010110010101100","0000111010001110100011101000","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000100100111001001110010011","0000100110011001100110011001","0000100000101000001010000010","0000011100000111000001110000","0000100110111001101110011011","0000010101100101011001010110","0001000000000000000000000000","0000101000011010000110100001","0000011110010111100101111001","0000100010101000101010001010","0000101000001010000010100000","0000100110111001101110011011","0000110010011100100111001001","0000100101111001011110010111","0000100000101000001010000010","0000101101011011010110110101","0000011001100110011001100110","0000010011110100111101001111","0000010110110101101101011011","0000100000111000001110000011","0000011100110111001101110011","0000000001010000010100000101","0000010110000101100001011000","0000111011111110111111101111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111111101111111011111110","0000101100111011001110110011","0000000110010001100100011001","0000000010100000101000001010","0001000000000000000000000000","0000000100100001001000010010","0000010010010100100101001001","0000100101111001011110010111","0000110010111100101111001011","0000110110001101100011011000","0000110101101101011011010110","0000110101111101011111010111","0000101110111011101110111011","0000100111111001111110011111","0000010001010100010101000101","0000001110000011100000111000","0000010101000101010001010100","0000010101010101010101010101","0000100010101000101010001010","0000100001001000010010000100","0000010110000101100001011000","0000011011010110110101101101","0000101000101010001010100010","0000110001001100010011000100","0000110111101101111011011110","0000111110101111101011111010","0000111011001110110011101100","0000110101001101010011010100","0000110001001100010011000100","0000110011001100110011001100","0000110110011101100111011001","0000110100101101001011010010","0000101111101011111010111110","0000101011001010110010101100","0000100101001001010010010100","0000101011011010110110101101","0000111100011111000111110001","0000111111111111111111111111","0000111100101111001011110010","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111101101111011011110110","0000110010111100101111001011","0000100110011001100110011001","0000101000011010000110100001","0000110010111100101111001011","0000110110111101101111011011","0000111100101111001011110010","0000110001011100010111000101","0000101100001011000010110000","0000011110100111101001111010","0000100111001001110010011100","0000100100101001001010010010","0000111010011110100111101001","0000111010101110101011101010","0000101110101011101010111010","0000110100101101001011010010","0000110011001100110011001100","0000111001111110011111100111","0000101011011010110110101101","0000101101101011011010110110","0000100110101001101010011010","0000011111100111111001111110","0000001001100010011000100110","0000001100010011000100110001","0000010101110101011101010111","0000000010010000100100001001","0000010001010100010101000101","0000011111000111110001111100","0000010100100101001001010010","0000011110010111100101111001","0000100001011000010110000101","0000100000001000000010000000","0000101101001011010010110100","0000110011001100110011001100","0000110110011101100111011001","0000110001011100010111000101","0000100011011000110110001101","0000101010001010100010101000","0000110100101101001011010010","0000111000011110000111100001","0000100110111001101110011011","0000010110110101101101011011","0000011001000110010001100100","0000111001011110010111100101","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111001111110011111100111","0000111110101111101011111010","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000110000011100000111000001","0000010011000100110001001100","0000000010000000100000001000","0000101010011010100110101001","0000111111011111110111111101","0000111111011111110111111101","0000111001101110011011100110","0000111011101110111011101110","0000111111111111111111111111","0000111010101110101011101010","0000101100011011000110110001","0000111100011111000111110001","0000111011111110111111101111","0000111111111111111111111111","0000111011001110110011101100","0000111100111111001111110011","0000111111011111110111111101","0000101010101010101010101010","0000011000000110000001100000","0000001010010010100100101001","0000010011010100110101001101","0000010111100101111001011110","0001000000000000000000000000","0000101001001010010010100100","0000100010111000101110001011","0000010110010101100101011001","0000110000011100000111000001","0000011011110110111101101111","0000011011110110111101101111","0000100000111000001110000011","0000011111100111111001111110","0000100111111001111110011111","0000011101000111010001110100","0000001001000010010000100100","0000001110100011101000111010","0000001011000010110000101100","0000000100100001001000010010","0001000000000000000000000000","0000010000000100000001000000","0000110011001100110011001100","0000111100001111000011110000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111011011110110111101101","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000110110001101100011011000","0000001010110010101100101011","0000000011000000110000001100","0001000000000000000000000000","0001000000000000000000000000","0000100000101000001010000010","0000110100101101001011010010","0000111110111111101111111011","0000111101001111010011110100","0000111010111110101111101011","0000111110111111101111111011","0000111101011111010111110101","0000110010001100100011001000","0000100100011001000110010001","0000011011010110110101101101","0000011111110111111101111111","0000011001010110010101100101","0000010010100100101001001010","0000011010010110100101101001","0000011110000111100001111000","0000110001001100010011000100","0000101111101011111010111110","0000101011111010111110101111","0000101010111010101110101011","0000110010101100101011001010","0000110110101101101011011010","0000110011101100111011001110","0000110001111100011111000111","0000110011001100110011001100","0000110001011100010111000101","0000101100111011001110110011","0000101001011010010110100101","0000111000001110000011100000","0000111111111111111111111111","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110101101101011011010","0000101100011011000110110001","0000101010101010101010101010","0000110101001101010011010100","0000110000101100001011000010","0000110110101101101011011010","0000111001101110011011100110","0000111010101110101011101010","0000101100101011001010110010","0000110111101101111011011110","0000100100011001000110010001","0000110011011100110111001101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100011111000111110001","0000110101001101010011010100","0000101110001011100010111000","0000101100011011000110110001","0000011010010110100101101001","0000011000000110000001100000","0000001111110011111100111111","0000001001110010011100100111","0001000000000000000000000000","0000001100000011000000110000","0000001100010011000100110001","0000010101110101011101010111","0000011000010110000101100001","0000011101110111011101110111","0000101101111011011110110111","0000101111101011111010111110","0000110011101100111011001110","0000111001101110011011100110","0000111101001111010011110100","0000111111111111111111111111","0000111011111110111111101111","0000101010111010101110101011","0000110000001100000011000000","0000111100111111001111110011","0000110101011101010111010101","0000100110111001101110011011","0000010010110100101101001011","0000100001111000011110000111","0000110110001101100011011000","0000111011111110111111101111","0000111111111111111111111111","0000111110001111100011111000","0000110111111101111111011111","0000110100101101001011010010","0000011011000110110001101100","0000000010100000101000001010","0000000100100001001000010010","0000101100111011001110110011","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111110101111101011111010","0000111010101110101011101010","0000111001111110011111100111","0000111010011110100111101001","0000110000001100000011000000","0000111001111110011111100111","0000111100001111000011110000","0000110110101101101011011010","0000111000011110000111100001","0000101010011010100110101001","0000011011110110111101101111","0000010000100100001001000010","0000001110010011100100111001","0000010011010100110101001101","0001000000000000000000000000","0000011111010111110101111101","0000100101011001010110010101","0000010110000101100001011000","0000101110001011100010111000","0000100100001001000010010000","0000010011110100111101001111","0000010101010101010101010101","0000011000010110000101100001","0000001100000011000000110000","0000001110100011101000111010","0000001100100011001000110010","0000001100010011000100110001","0000001010010010100100101001","0000000110000001100000011000","0000000011000000110000001100","0000011111010111110101111101","0000111111111111111111111111","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111011101110111011101110","0000111101011111010111110101","0000111111111111111111111111","0000111011111110111111101111","0000011101100111011001110110","0000000101000001010000010100","0001000000000000000000000000","0001000000000000000000000000","0000100110111001101110011011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111001111110011111100","0000111011001110110011101100","0000111111111111111111111111","0000110101111101011111010111","0000100010111000101110001011","0000011110000111100001111000","0000010111000101110001011100","0001000000000000000000000000","0000100111001001110010011100","0000101101101011011010110110","0000110000111100001111000011","0000110000111100001111000011","0000110111101101111011011110","0000110000101100001011000010","0000101010001010100010101000","0000101001101010011010100110","0000101100111011001110110011","0000101111111011111110111111","0000110000101100001011000010","0000110000111100001111000011","0000111110001111100011111000","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111110111111101111111011","0000111100111111001111110011","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000101011101010111010101110","0000101101001011010010110100","0000111111111111111111111111","0000110010001100100011001000","0000111101001111010011110100","0000111110101111101011111010","0000111000111110001111100011","0000111100101111001011110010","0000110100001101000011010000","0000110110101101101011011010","0000110101101101011011010110","0000110000001100000011000000","0000110111111101111111011111","0000111010101110101011101010","0000111010011110100111101001","0000111111111111111111111111","0000111111001111110011111100","0000101101011011010110110101","0000101010101010101010101010","0000011000000110000001100000","0000100100111001001110010011","0000001011000010110000101100","0000001010100010101000101010","0000001101000011010000110100","0000001101110011011100110111","0000000111110001111100011111","0000001001100010011000100110","0000011000000110000001100000","0000100000001000000010000000","0000101100101011001010110010","0000111101101111011011110110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000110100011101000111010001","0000111000001110000011100000","0000110101101101011011010110","0000110101001101010011010100","0000011100010111000101110001","0000001000110010001100100011","0000001110000011100000111000","0000010001000100010001000100","0000010011000100110001001100","0000001110100011101000111010","0000000011000000110000001100","0000000000110000001100000011","0000010110110101101101011011","0000110011111100111111001111","0000110101101101011011010110","0000111101011111010111110101","0000111011011110110111101101","0000111110101111101011111010","0000111101011111010111110101","0000111111111111111111111111","0000111101001111010011110100","0000111100111111001111110011","0000110010111100101111001011","0000110000111100001111000011","0000110000111100001111000011","0000101110001011100010111000","0000110000011100000111000001","0000100100001001000010010000","0000100111101001111010011110","0000011011110110111101101111","0000001110010011100100111001","0000001011000010110000101100","0000000100110001001100010011","0000011011010110110101101101","0000100101001001010010010100","0000101011101010111010101110","0000010010110100101101001011","0000101000101010001010100010","0000011100000111000001110000","0000010011100100111001001110","0000000011110000111100001111","0000000011010000110100001101","0000011010110110101101101011","0000001101000011010000110100","0000101000011010000110100001","0000001011100010111000101110","0001000000000000000000000000","0000000111010001110100011101","0000101110101011101010111010","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111100111111001111110011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111111001111110011111100","0000111110011111100111111001","0000111100011111000111110001","0000111011111110111111101111","0000111100111111001111110011","0000111100011111000111110001","0000111111111111111111111111","0000111101001111010011110100","0000111110001111100011111000","0000101010101010101010101010","0001000000000000000000000000","0000000010110000101100001011","0000000010010000100100001001","0000101100111011001110110011","0000111111111111111111111111","0000111101111111011111110111","0000111001001110010011100100","0000111111111111111111111111","0000111101011111010111110101","0000111110101111101011111010","0000111111001111110011111100","0000111000011110000111100001","0000100101101001011010010110","0000101100011011000110110001","0000000101000001010000010100","0000101011111010111110101111","0000101100011011000110110001","0000111010101110101011101010","0000110101001101010011010100","0000101011001010110010101100","0000110100101101001011010010","0000111001101110011011100110","0000110001011100010111000101","0000100101101001011010010110","0000100110001001100010011000","0000110100011101000111010001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111001111110011111100","0000111111101111111011111110","0000111111011111110111111101","0000111110011111100111111001","0000111111011111110111111101","0000111111001111110011111100","0000111111001111110011111100","0000111110101111101011111010","0000110110101101101011011010","0000101000111010001110100011","0000111111111111111111111111","0000111001011110010111100101","0000110110101101101011011010","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111011011110110111101101","0000111011001110110011101100","0000110100001101000011010000","0000111010001110100011101000","0000110011111100111111001111","0000110011101100111011001110","0000101000011010000110100001","0000110110101101101011011010","0000111101001111010011110100","0000110110011101100111011001","0000100011001000110010001100","0000001010000010100000101000","0000011001110110011101100111","0000010001100100011001000110","0000001101100011011000110110","0000010101110101011101010111","0000010001100100011001000110","0000001111100011111000111110","0000010001100100011001000110","0000011111010111110101111101","0000101010101010101010101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111011101110111011101110","0000111111111111111111111111","0000111100011111000111110001","0000111100001111000011110000","0000111100011111000111110001","0000111111111111111111111111","0000111001001110010011100100","0000110111101101111011011110","0000101101111011011110110111","0000101101101011011010110110","0000101010111010101110101011","0000011100110111001101110011","0000011101000111010001110100","0000010110110101101101011011","0000010000100100001001000010","0000011001000110010001100100","0000101011111010111110101111","0000110100001101000011010000","0000110000101100001011000010","0000111010111110101111101011","0000111111101111111011111110","0000111111111111111111111111","0000111110001111100011111000","0000111101011111010111110101","0000111111111111111111111111","0000101101001011010010110100","0000101011101010111010101110","0000100001101000011010000110","0000011100010111000101110001","0000011111100111111001111110","0000011111100111111001111110","0000011100000111000001110000","0000101010101010101010101010","0000011110000111100001111000","0000001110100011101000111010","0000000101000001010000010100","0000001010100010101000101010","0000011001110110011101100111","0000101011111010111110101111","0000100010111000101110001011","0000010000100100001001000010","0000101110101011101010111010","0000010010110100101101001011","0000011100000111000001110000","0000001000010010000100100001","0000001111100011111000111110","0000100111011001110110011101","0000110010111100101111001011","0000001100000011000000110000","0001000000000000000000000000","0000000000100000001000000010","0000001101110011011100110111","0000110000001100000011000000","0000111100101111001011110010","0000111111111111111111111111","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111011111110111111101","0000111111111111111111111111","0000111101011111010111110101","0000111100011111000111110001","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000110001001100010011000100","0001000000000000000000000000","0000000011010000110100001101","0000001001010010010100100101","0000110100011101000111010001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000101101111011011110110111","0000001010000010100000101000","0000100110101001101010011010","0000110110101101101011011010","0000111000111110001111100011","0000111111111111111111111111","0000111010111110101111101011","0000110111001101110011011100","0000101110111011101110111011","0000101010011010100110101001","0000110001111100011111000111","0000111110101111101011111010","0000111111111111111111111111","0000111110011111100111111001","0000111100111111001111110011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111110001111100011111000","0000111011111110111111101111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111011011110110111101101","0000101100111011001110110011","0000101111001011110010111100","0000101111001011110010111100","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111001111110011111100111","0000111011001110110011101100","0000111100101111001011110010","0000111110001111100011111000","0000110010101100101011001010","0000111111111111111111111111","0000110101001101010011010100","0000101000101010001010100010","0000011000010110000101100001","0000000111010001110100011101","0000011100100111001001110010","0001000000000000000000000000","0000001000110010001100100011","0000001001110010011100100111","0000000110100001101000011010","0000010001110100011101000111","0000010100110101001101010011","0000110100111101001111010011","0000111100111111001111110011","0000111111111111111111111111","0000111101101111011011110110","0000111110011111100111111001","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011101110111011101110","0000111111111111111111111111","0000111111101111111011111110","0000110110001101100011011000","0000100011101000111010001110","0000011010010110100101101001","0000100101011001010110010101","0000100111011001110110011101","0000100011011000110110001101","0000011101110111011101110111","0000100001101000011010000110","0000101100101011001010110010","0000111000001110000011100000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000101011101010111010101110","0000011010110110101101101011","0000011101110111011101110111","0000001110110011101100111011","0000011110010111100101111001","0000110100111101001111010011","0000101001101010011010100110","0000100011011000110110001101","0000000011000000110000001100","0001000000000000000000000000","0000000100100001001000010010","0000011010110110101101101011","0000011010110110101101101011","0000100010001000100010001000","0000100001001000010010000100","0000100011011000110110001101","0000100100101001001010010010","0000011110100111101001111010","0000011101010111010101110101","0000011011100110111001101110","0000011000110110001101100011","0000011100100111001001110010","0000100000011000000110000001","0000100100101001001010010010","0000010010100100101001001010","0000011000000110000001100000","0001000000000000000000000000","0000100100101001001010010010","0000101110111011101110111011","0000111100111111001111110011","0000111111111111111111111111","0000111101111111011111110111","0000111101101111011011110110","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111011101110111011101110","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110001111100011111000","0000111111001111110011111100","0000111111111111111111111111","0000111011111110111111101111","0000111101011111010111110101","0000111110001111100011111000","0000111110011111100111111001","0000110110111101101111011011","0000000110010001100100011001","0001000000000000000000000000","0001000000000000000000000000","0000100000111000001110000011","0000111010101110101011101010","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111101011111010111110101","0000111111111111111111111111","0000110110101101101011011010","0000110010111100101111001011","0000010010100100101001001010","0000011001110110011101100111","0000111111111111111111111111","0000111100111111001111110011","0000111110101111101011111010","0000110111111101111111011111","0000111001011110010111100101","0000111011101110111011101110","0000111101101111011011110110","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111110101111101011111010","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111111101111111011111110","0000111111001111110011111100","0000111100101111001011110010","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111101011111010111110101","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000110110101101101011011010","0000101001011010010110100101","0000110110001101100011011000","0000110100001101000011010000","0000110010001100100011001000","0000110111101101111011011110","0000111101011111010111110101","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000110101101101011011010110","0000111100101111001011110010","0000110101101101011011010110","0000011101100111011001110110","0000011100010111000101110001","0000001011100010111000101110","0000100110011001100110011001","0001000000000000000000000000","0000001000110010001100100011","0000010011100100111001001110","0000001011000010110000101100","0000010010100100101001001010","0000011001100110011001100110","0000111110101111101011111010","0000111111111111111111111111","0000111100001111000011110000","0000111111001111110011111100","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111111001111110011111100","0000111110111111101111111011","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000110000111100001111000011","0000101010011010100110101001","0000110000001100000011000000","0000111010011110100111101001","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000110010001100100011001000","0000011011000110110001101100","0000010110010101100101011001","0000010001010100010101000101","0000001011010010110100101101","0000011101100111011001110110","0000101011001010110010101100","0000100011001000110010001100","0000101001101010011010100110","0000101111001011110010111100","0000110001011100010111000101","0000111100111111001111110011","0000111111001111110011111100","0000100001111000011110000111","0000100100101001001010010010","0000101100111011001110110011","0000101101001011010010110100","0000011001000110010001100100","0000110001111100011111000111","0000010110100101101001011010","0000011011100110111001101110","0000001111110011111100111111","0000010110100101101001011010","0000011111010111110101111101","0000010011110100111101001111","0000000001110000011100000111","0000011100010111000101110001","0000000011110000111100001111","0000101100011011000110110001","0000111010101110101011101010","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111001111110011111100","0000111110101111101011111010","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000010110100101101001011010","0000000001110000011100000111","0001000000000000000000000000","0000001100000011000000110000","0000101110011011100110111001","0000111111111111111111111111","0000111011111110111111101111","0000111110101111101011111010","0000111101101111011011110110","0000111100101111001011110010","0000101111111011111110111111","0000010100000101000001010000","0000100000011000000110000001","0000111111011111110111111101","0000111101101111011011110110","0000110110111101101111011011","0000101100111011001110110011","0000111100011111000111110001","0000111110001111100011111000","0000111101111111011111110111","0000110101101101011011010110","0000110110101101101011011010","0000110001101100011011000110","0000110110111101101111011011","0000110111111101111111011111","0000111000111110001111100011","0000111010111110101111101011","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111110111111101111111011","0000111100101111001011110010","0000110110111101101111011011","0000101101101011011010110110","0000101011001010110010101100","0000100011011000110110001101","0000011100000111000001110000","0000010011110100111101001111","0000011001110110011101100111","0000100000111000001110000011","0000100101011001010110010101","0000100101101001011010010110","0000110100001101000011010000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111001011110010111100101","0000111001101110011011100110","0000101001111010011110100111","0000100011011000110110001101","0000010011000100110001001100","0000010001000100010001000100","0000000111100001111000011110","0000100100011001000110010001","0001000000000000000000000000","0000000001000000010000000100","0000011111000111110001111100","0000011011010110110101101101","0000010110010101100101011001","0000001111000011110000111100","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101001111010011110100","0000111110011111100111111001","0000111010001110100011101000","0000111111111111111111111111","0000111110001111100011111000","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111100101111001011110010","0000111101111111011111110111","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111100001111000011110000","0000111101111111011111110111","0000111111101111111011111110","0000111101101111011011110110","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111100001111000011110000","0000101100111011001110110011","0000010110010101100101011001","0000001101100011011000110110","0000011000010110000101100001","0000100110111001101110011011","0000110100001101000011010000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000111100111111001111110011","0000111111111111111111111111","0000101101111011011110110111","0000011111110111111101111111","0000111100111111001111110011","0000101000101010001010100010","0000011110000111100001111000","0000101101111011011110110111","0000100011101000111010001110","0000001011000010110000101100","0000100001111000011110000111","0000010110000101100001011000","0000010010110100101101001011","0000101000101010001010100010","0001000000000000000000000000","0000000010000000100000001000","0000110010011100100111001001","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000101010111010101110101011","0000011001100110011001100110","0000000111010001110100011101","0000000000010000000100000001","0000011001110110011101100111","0000110101001101010011010100","0000111001001110010011100100","0000111110101111101011111010","0000111011101110111011101110","0000101011101010111010101110","0000011000100110001001100010","0000010010100100101001001010","0000110010011100100111001001","0000110111011101110111011101","0000101100101011001010110010","0000100101011001010110010101","0000100111001001110010011100","0000100110111001101110011011","0000100101101001011010010110","0000101000001010000010100000","0000100110101001101010011010","0000011111100111111001111110","0000010111100101111001011110","0000010101110101011101010111","0000011010110110101101101011","0000100001001000010010000100","0000100101101001011010010110","0000101000001010000010100000","0000101010111010101110101011","0000101110101011101010111010","0000110001101100011011000110","0000110000101100001011000010","0000110100101101001011010010","0000110111011101110111011101","0000110001011100010111000101","0000110110001101100011011000","0000101101111011011110110111","0000011110100111101001111010","0000011011110110111101101111","0000010100010101000101010001","0000001001010010010100100101","0000001011110010111100101111","0000100010001000100010001000","0000011110000111100001111000","0000100100101001001010010010","0000100101001001010010010100","0000100110111001101110011011","0000110110011101100111011001","0000101010101010101010101010","0000100011011000110110001101","0000011111010111110101111101","0000010011000100110001001100","0000100011111000111110001111","0000011010000110100001101000","0000001000110010001100100011","0000010001100100011001000110","0000101011111010111110101111","0001000000000000000000000000","0000001000000010000000100000","0000010110000101100001011000","0000010101110101011101010111","0000101000101010001010100010","0000001110100011101000111010","0000110101011101010111010101","0000111111111111111111111111","0000111111001111110011111100","0000111010011110100111101001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111111001111110011111100","0000111101111111011111110111","0000111111111111111111111111","0000111011011110110111101101","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101001111010011110100","0000111111111111111111111111","0000111001011110010111100101","0000111101001111010011110100","0000111101101111011011110110","0000111101011111010111110101","0000101100011011000110110001","0000010000000100000001000000","0000010000110100001101000011","0000100110111001101110011011","0000110010011100100111001001","0000111101001111010011110100","0000111111111111111111111111","0000111010111110101111101011","0000111110111111101111111011","0000111010111110101111101011","0000111011011110110111101101","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111100111111001111110011","0000110110101101101011011010","0000100100101001001010010010","0000111110101111101011111010","0000101011101010111010101110","0000100100001001000010010000","0000110001111100011111000111","0000011100000111000001110000","0000010101010101010101010101","0000011110010111100101111001","0000010101110101011101010111","0000100001011000010110000101","0000011001100110011001100110","0000000001110000011100000111","0000101100001011000010110000","0000111101001111010011110100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000110010011100100111001001","0000011000110110001101100011","0000010010110100101101001011","0000001101000011010000110100","0000000011110000111100001111","0000010011010100110101001101","0000011110110111101101111011","0000101001101010011010100110","0000100100111001001110010011","0000001000000010000000100000","0000101000111010001110100011","0000110110011101100111011001","0000011100010111000101110001","0000010101110101011101010111","0000011101100111011001110110","0000100011001000110010001100","0000100011101000111010001110","0000010111110101111101011111","0000001100100011001000110010","0000001000000010000000100000","0000001001100010011000100110","0000001000110010001100100011","0001000000000000000000000000","0001000000000000000000000000","0000000010010000100100001001","0000001001000010010000100100","0000010000110100001101000011","0000010110000101100001011000","0000010111000101110001011100","0000010110010101100101011001","0000011101000111010001110100","0000100110111001101110011011","0000100111111001111110011111","0000101111001011110010111100","0000011010000110100001101000","0000100100001001000010010000","0000100101101001011010010110","0000010100010101000101010001","0000010000100100001001000010","0000010100010101000101010001","0000001101100011011000110110","0000010001000100010001000100","0000101110111011101110111011","0000110001101100011011000110","0000101000011010000110100001","0000101001011010010110100101","0000011011100110111001101110","0000011111100111111001111110","0000100010111000101110001011","0000001100100011001000110010","0000010111000101110001011100","0000010000010100000101000001","0000010010010100100101001001","0000100100101001001010010010","0000100001111000011110000111","0000111010101110101011101010","0000000010010000100100001001","0000100100001001000010010000","0000000101110001011100010111","0001000000000000000000000000","0000100110011001100110011001","0000100111111001111110011111","0000100110011001100110011001","0000111111111111111111111111","0000111101001111010011110100","0000110101011101010111010101","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111100001111000011110000","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000110111111101111111011111","0000111101001111010011110100","0000111111111111111111111111","0000111100101111001011110010","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000101011101010111010101110","0000010001010100010101000101","0000011010110110101101101011","0000101100101011001010110010","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111011001110110011101100","0000111111111111111111111111","0000111011101110111011101110","0000111111111111111111111111","0000111000111110001111100011","0000101010011010100110101001","0000110100101101001011010010","0000111101111111011111110111","0000110000011100000111000001","0000100111001001110010011100","0000101001001010010010100100","0000100011001000110010001100","0000011001010110010101100101","0000100111001001110010011100","0000011000100110001001100010","0000100001011000010110000101","0000000000100000001000000010","0000101011001010110010101100","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110001111100011111000","0000111100101111001011110010","0000111111111111111111111111","0000100110101001101010011010","0000001100000011000000110000","0000001100000011000000110000","0001000000000000000000000000","0000001100100011001000110010","0000011101010111010101110101","0000100000101000001010000010","0000000110100001101000011010","0000010000100100001001000010","0000000100110001001100010011","0000000111100001111000011110","0000001010000010100000101000","0001000000000000000000000000","0000000010010000100100001001","0000000011100000111000001110","0000000111010001110100011101","0000011001000110010001100100","0000100111111001111110011111","0000100111101001111010011110","0000011111010111110101111101","0000110001101100011011000110","0000110011111100111111001111","0000110110111101101111011011","0000111001001110010011100100","0000111010101110101011101010","0000111011101110111011101110","0000111101001111010011110100","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111010011110100111101001","0000101111001011110010111100","0000110111011101110111011101","0000101000011010000110100001","0000011101100111011001110110","0000110101111101011111010111","0000111000001110000011100000","0000100011001000110010001100","0000010011100100111001001110","0000011110100111101001111010","0000001110100011101000111010","0000101001111010011110100111","0000101111001011110010111100","0000100110101001101010011010","0000011110000111100001111000","0000010101100101011001010110","0000100010101000101010001010","0000011100010111000101110001","0000010111100101111001011110","0000100000001000000010000000","0000101010011010100110101001","0000011111010111110101111101","0000100100001001000010010000","0000101101001011010010110100","0000000001000000010000000100","0000100111011001110110011101","0000010010010100100101001001","0000001101110011011100110111","0000010100110101001101010011","0000110111111101111111011111","0000100100001001000010010000","0000110011011100110111001101","0000111011001110110011101100","0000110011011100110111001101","0000111011101110111011101110","0000111100111111001111110011","0000111111111111111111111111","0000111101001111010011110100","0000110101111101011111010111","0000110000011100000111000001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111011011110110111101101","0000111111111111111111111111","0000110010001100100011001000","0000010011010100110101001101","0000011010110110101101101011","0000111001101110011011100110","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111011111110111111101","0000111000111110001111100011","0000111111111111111111111111","0000111111111111111111111111","0000111100101111001011110010","0000111110011111100111111001","0000111111111111111111111111","0000111101011111010111110101","0000111000101110001011100010","0000111000111110001111100011","0000101010111010101110101011","0000111111111111111111111111","0000111101001111010011110100","0000110100011101000111010001","0000100110001001100010011000","0000101011001010110010101100","0000101100011011000110110001","0000011111110111111101111111","0000101101011011010110110101","0000011100110111001101110011","0000000111000001110000011100","0000011111100111111001111110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111110011111100111111001","0000111110011111100111111001","0000111111001111110011111100","0000111111111111111111111111","0000111010001110100011101000","0000100110101001101010011010","0000011011110110111101101111","0000001101000011010000110100","0001000000000000000000000000","0001000000000000000000000000","0000000011010000110100001101","0000001011100010111000101110","0000010111100101111001011110","0001000000000000000000000000","0000000001100000011000000110","0000010111110101111101011111","0000101000011010000110100001","0000110100011101000111010001","0000100000011000000110000001","0000101011001010110010101100","0000100111111001111110011111","0000110110101101101011011010","0000111001111110011111100111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000110001011100010111000101","0000111000001110000011100000","0000110111011101110111011101","0000111001101110011011100110","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111010111110101111101011","0000110000001100000011000000","0001000000000000000000000000","0000000011100000111000001110","0000011001010110010101100101","0000111111111111111111111111","0000111001111110011111100111","0000110011001100110011001100","0000101001011010010110100101","0000110001111100011111000111","0000100011101000111010001110","0000101110011011100110111001","0000011110000111100001111000","0000100110011001100110011001","0000001110110011101100111011","0000100011011000110110001101","0000011000000110000001100000","0000001110100011101000111010","0000010000110100001101000011","0000010010110100101101001011","0000100010011000100110001001","0000010001100100011001000110","0000100010111000101110001011","0000101101011011010110110101","0000101011111010111110101111","0000101100111011001110110011","0000101001001010010010100100","0000111111111111111111111111","0000111001001110010011100100","0000110110011101100111011001","0000110111011101110111011101","0000101111111011111110111111","0000111110001111100011111000","0000111101011111010111110101","0000111110011111100111111001","0000111111111111111111111111","0000111100001111000011110000","0000111110011111100111111001","0000111111111111111111111111","0000110111101101111011011110","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000110111101101111011011110","0000011011010110110101101101","0000001101010011010100110101","0000111001101110011011100110","0000111111011111110111111101","0000111110101111101011111010","0000111100001111000011110000","0000111111001111110011111100","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111010011110100111101001","0000111110001111100011111000","0000111001101110011011100110","0000111000111110001111100011","0000110010101100101011001010","0000111100101111001011110010","0000101011011010110110101101","0000111111111111111111111111","0000111110101111101011111010","0000110110111101101111011011","0000100100001001000010010000","0000111110011111100111111001","0000101101111011011110110111","0000101010001010100010101000","0000100101001001010010010100","0000001111000011110000111100","0000010111010101110101011101","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000111111111111111111111111","0000111100111111001111110011","0000111110011111100111111001","0000111110111111101111111011","0000111011011110110111101101","0000111111111111111111111111","0000111110011111100111111001","0000111111101111111011111110","0000111110011111100111111001","0000101101001011010010110100","0000000000010000000100000001","0000010010100100101001001010","0000000101100001011000010110","0000010011010100110101001101","0000100011111000111110001111","0000100000111000001110000011","0000100110101001101010011010","0000011100110111001101110011","0000100100101001001010010010","0000101100001011000010110000","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111100111111001111110011","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111110011111100111111001","0000111011111110111111101111","0000111111001111110011111100","0000101001101010011010100110","0000111001101110011011100110","0000111010111110101111101011","0000111110001111100011111000","0000111010001110100011101000","0000111111111111111111111111","0000111101001111010011110100","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000100011101000111010001110","0000011110100111101001111010","0000010101010101010101010101","0000101101111011011110110111","0000111110101111101011111010","0000111111111111111111111111","0000111110111111101111111011","0000111110011111100111111001","0000111001101110011011100110","0000101001101010011010100110","0000010111000101110001011100","0000011010110110101101101011","0000001101100011011000110110","0000100101011001010110010101","0000010001110100011101000111","0000100001101000011010000110","0000100001011000010110000101","0001000000000000000000000000","0000001011100010111000101110","0000100000101000001010000010","0000000000110000001100000011","0000010110100101101001011010","0000011001000110010001100100","0000101101101011011010110110","0000101001001010010010100100","0000101110111011101110111011","0000110011011100110111001101","0000111101111111011111110111","0000110010111100101111001011","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111110101111101011111010","0000110010111100101111001011","0000111111111111111111111111","0000111000011110000111100001","0000111000101110001011100010","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000111001001110010011100100","0000111111111111111111111111","0000010101100101011001010110","0000001101110011011100110111","0000111000111110001111100011","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101101111011011110110","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111001111110011111100111","0000110000011100000111000001","0000111111111111111111111111","0000100011101000111010001110","0000111010111110101111101011","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111010001110100011101000","0000100100011001000110010001","0000111111101111111011111110","0000110110101101101011011010","0000100011111000111110001111","0000011100010111000101110001","0000000111110001111100011111","0000111100001111000011110000","0000111110011111100111111001","0000111111111111111111111111","0000111101111111011111110111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111111101111111011111110","0000111111111111111111111111","0000111101101111011011110110","0000111101111111011111110111","0000111011111110111111101111","0000111001011110010111100101","0000111011001110110011101100","0000111111111111111111111111","0000111110111111101111111011","0000011110100111101001111010","0001000000000000000000000000","0000010010110100101101001011","0000010101010101010101010101","0000011101000111010001110100","0000011111110111111101111111","0000010101010101010101010101","0000100000101000001010000010","0000101100111011001110110011","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111001101110011011100110","0000111100111111001111110011","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000110011111100111111001111","0000111110001111100011111000","0000111111011111110111111101","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111110001111100011111000","0000111111111111111111111111","0000111110111111101111111011","0000111011101110111011101110","0000100001001000010010000100","0000011110010111100101111001","0000100100101001001010010010","0000110110111101101111011011","0000111000111110001111100011","0000111110111111101111111011","0000111110101111101011111010","0000101100011011000110110001","0000101000101010001010100010","0000100111111001111110011111","0000101010011010100110101001","0000001111100011111000111110","0000100010011000100110001001","0000001001100010011000100110","0000100101101001011010010110","0000111111111111111111111111","0000010000100100001001000010","0000000001100000011000000110","0000100000111000001110000011","0001000000000000000000000000","0000010110000101100001011000","0000000011110000111100001111","0000001000100010001000100010","0000011011010110110101101101","0000101011101010111010101110","0000101010001010100010101000","0000101100101011001010110010","0000111001101110011011100110","0000111010001110100011101000","0000111001111110011111100111","0000111011001110110011101100","0000110101011101010111010101","0000110010001100100011001000","0000111010011110100111101001","0000110011011100110111001101","0000111111001111110011111100","0000111111111111111111111111","0000110000111100001111000011","0000110111011101110111011101","0000110000101100001011000010","0000000011100000111000001110","0000010110110101101101011011","0000111101001111010011110100","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111100101111001011110010","0000111001001110010011100100","0000100011001000110010001100","0000111000011110000111100001","0000101110011011100110111001","0000011100100111001001110010","0000011100110111001101110011","0000100111011001110110011101","0000111101011111010111110101","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000101001001010010010100100","0000110101111101011111010111","0000111101001111010011110100","0000010110000101100001011000","0000001111110011111100111111","0000100001011000010110000101","0000111101011111010111110101","0000111101111111011111110111","0000111111011111110111111101","0000111100101111001011110010","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111100111111001111110011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111011101110111011101110","0001000000000000000000000000","0000011000000110000001100000","0000011101000111010001110100","0000010011100100111001001110","0000011000100110001001100010","0000001011100010111000101110","0000011000010110000101100001","0000111101011111010111110101","0000111100011111000111110001","0000111111111111111111111111","0000111100001111000011110000","0000110111011101110111011101","0000111111111111111111111111","0000111111101111111011111110","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111001001110010011100100","0000111111111111111111111111","0000111111001111110011111100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111011101110111011101110","0000111111111111111111111111","0000101010111010101110101011","0000100100011001000110010001","0000100001011000010110000101","0000100110101001101010011010","0000101001111010011110100111","0000111110111111101111111011","0000111010111110101111101011","0000101001101010011010100110","0000100100111001001110010011","0000101010001010100010101000","0000100010111000101110001011","0000011101010111010101110101","0000100100011001000110010001","0000000101100001011000010110","0000101100111011001110110011","0000111110101111101011111010","0000111010001110100011101000","0000001101010011010100110101","0000001001010010010100100101","0000011110100111101001111010","0000011110000111100001111000","0000010101100101011001010110","0000001101000011010000110100","0000000110010001100100011001","0000000001000000010000000100","0000010100000101000001010000","0000100000001000000010000000","0000101100011011000110110001","0000110101011101010111010101","0000110110111101101111011011","0000100111001001110010011100","0000110001011100010111000101","0000111011001110110011101100","0000101011111010111110101111","0000111111111111111111111111","0000110001101100011011000110","0000011111110111111101111111","0000100001001000010010000100","0000001010110010101100101011","0000000100100001001000010010","0000101011101010111010101110","0000111100101111001011110010","0000111001111110011111100111","0000111111101111111011111110","0000111111111111111111111111","0000111100101111001011110010","0000111101101111011011110110","0000111111001111110011111100","0000111101101111011011110110","0000111110111111101111111011","0000111111111111111111111111","0000111101111111011111110111","0000100011011000110110001101","0000010101000101010001010100","0000110111001101110011011100","0000010111010101110101011101","0000011100000111000001110000","0000111101101111011011110110","0000111111111111111111111111","0000111100101111001011110010","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000110000001100000011000000","0000111001001110010011100100","0000110101001101010011010100","0000010011110100111101001111","0001000000000000000000000000","0000111000111110001111100011","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000111111101111111011111110","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111100111111001111110011","0000111101111111011111110111","0000111110101111101011111010","0000111110111111101111111011","0000101110011011100110111001","0000000011010000110100001101","0000001011000010110000101100","0000011010010110100101101001","0000010100100101001001010010","0000010010100100101001001010","0000011000110110001101100011","0000101111001011110010111100","0000111110111111101111111011","0000111110101111101011111010","0000110111101101111011011110","0000111010011110100111101001","0000111011001110110011101100","0000111111111111111111111111","0000111101101111011011110110","0000111011001110110011101100","0000111111001111110011111100","0000111010101110101011101010","0000111111011111110111111101","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111011111110111111101","0000111110111111101111111011","0000111101011111010111110101","0000111100101111001011110010","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111101101111011011110110","0000110111111101111111011111","0000100100011001000110010001","0000001110100011101000111010","0000011111110111111101111111","0000100111011001110110011101","0000101111111011111110111111","0000110010001100100011001000","0000110011011100110111001101","0000001010000010100000101000","0000011011110110111101101111","0000100011001000110010001100","0000100001111000011110000111","0000100111001001110010011100","0000000100010001000100010001","0000111001011110010111100101","0000111111001111110011111100","0000111111111111111111111111","0000111000001110000011100000","0000010011010100110101001101","0000001000000010000000100000","0001000000000000000000000000","0000010001110100011101000111","0000010001010100010101000101","0000001100010011000100110001","0000010100100101001001010010","0000001100100011001000110010","0001000000000000000000000000","0000000010000000100000001000","0000001101000011010000110100","0000010000100100001001000010","0000010100010101000101010001","0000010110100101101001011010","0000010001000100010001000100","0000011001100110011001100110","0000001101000011010000110100","0000000000110000001100000011","0001000000000000000000000000","0000010001110100011101000111","0000101001101010011010100110","0000111010101110101011101010","0000111111111111111111111111","0000111011111110111111101111","0000111000111110001111100011","0000111101001111010011110100","0000111111001111110011111100","0000111111111111111111111111","0000111101101111011011110110","0000111111101111111011111110","0000111110001111100011111000","0000111110111111101111111011","0000111010101110101011101010","0000100100101001001010010010","0000110001101100011011000110","0000010011000100110001001100","0000101100101011001010110010","0000001111110011111100111111","0000110110001101100011011000","0000111111111111111111111111","0000111110001111100011111000","0000111110001111100011111000","0000111101111111011111110111","0000111111011111110111111101","0000111110111111101111111011","0000111010001110100011101000","0000111010001110100011101000","0000011101110111011101110111","0001000000000000000000000000","0000011100100111001001110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111011101110111011101110","0000011011100110111001101110","0001000000000000000000000000","0000011010010110100101101001","0000011110110111101101111011","0000011011110110111101101111","0000100001001000010010000100","0000101010011010100110101001","0000101011101010111010101110","0000111111111111111111111111","0000111111111111111111111111","0000101110101011101010111010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000110111011101110111011101","0000111001101110011011100110","0000111100011111000111110001","0000111111111111111111111111","0000111110101111101011111010","0000111101111111011111110111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111100111111001111110011","0000111111111111111111111111","0000111011101110111011101110","0000110110001101100011011000","0000100110001001100010011000","0000001100100011001000110010","0000000010110000101100001011","0000000111000001110000011100","0000010000010100000101000001","0000011010000110100001101000","0000101011101010111010101110","0000101110001011100010111000","0000001001110010011100100111","0000000110100001101000011010","0000010100010101000101010001","0000011110000111100001111000","0000011110000111100001111000","0001000000000000000000000000","0000111111011111110111111101","0000111111111111111111111111","0000111000101110001011100010","0000111111111111111111111111","0000111101001111010011110100","0000010000110100001101000011","0000000001010000010100000101","0000010110010101100101011001","0000010010000100100001001000","0000010000010100000101000001","0000010000000100000001000000","0000001100000011000000110000","0000001010100010101000101010","0000001001000010010000100100","0000001001000010010000100100","0000000011100000111000001110","0000000001000000010000000100","0001000000000000000000000000","0000000111000001110000011100","0000001100010011000100110001","0000010001110100011101000111","0000101000101010001010100010","0000111000101110001011100010","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111100011111000111110001","0000111111111111111111111111","0000111011001110110011101100","0000110110111101101111011011","0000111110111111101111111011","0000111110111111101111111011","0000111111111111111111111111","0000111110101111101011111010","0000111110011111100111111001","0000110111001101110011011100","0000101111011011110110111101","0000111011001110110011101100","0000100101111001011110010111","0000001110010011100100111001","0000100011011000110110001101","0000001010110010101100101011","0000111000001110000011100000","0000101100101011001010110010","0000111101111111011111110111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110110011101100111011001","0000101110111011101110111011","0000011100110111001101110011","0000000001110000011100000111","0000100101111001011110010111","0000101100111011001110110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000110111111101111111011111","0000001100000011000000110000","0000000010110000101100001011","0000011100110111001101110011","0000011100000111000001110000","0000011011100110111001101110","0000101100011011000110110001","0000101100001011000010110000","0000110010011100100111001001","0000101111101011111010111110","0000110110111101101111011011","0000111100111111001111110011","0000111110111111101111111011","0000111100101111001011110010","0000111010101110101011101010","0000111110001111100011111000","0000101111011011110110111101","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111101111111011111110111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101001111010011110100","0000110000111100001111000011","0000101100111011001110110011","0000100111101001111010011110","0000010011100100111001001110","0000001011100010111000101110","0000000100000001000000010000","0000000100100001001000010010","0000000011110000111100001111","0001000000000000000000000000","0001000000000000000000000000","0000011110110111101101111011","0000001101000011010000110100","0000010001010100010101000101","0000001101110011011100110111","0000100000111000001110000011","0000000111110001111100011111","0000010110000101100001011000","0000111111111111111111111111","0000111100001111000011110000","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000110000011100000111000001","0001000000000000000000000000","0000000010100000101000001010","0000001001100010011000100110","0000010010010100100101001001","0000010001010100010101000101","0000010100110101001101010011","0000100000001000000010000000","0000100000101000001010000010","0000101111111011111110111111","0000011011010110110101101101","0000100001001000010010000100","0000100001101000011010000110","0000110101011101010111010101","0000111101101111011011110110","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111001101110011011100110","0000111111111111111111111111","0000111010101110101011101010","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111101011111010111110101","0000101111001011110010111100","0000110010001100100011001000","0000111010111110101111101011","0000110010111100101111001011","0000101110011011100110111001","0000111001111110011111100111","0000111000001110000011100000","0000101110001011100010111000","0000100011101000111010001110","0000011011110110111101101111","0000001111110011111100111111","0001000000000000000000000000","0000011000110110001101100011","0000111110011111100111111001","0000111110111111101111111011","0000111010111110101111101011","0000101111101011111010111110","0000101110111011101110111011","0000011101100111011001110110","0000100001111000011110000111","0000100100101001001010010010","0000010001110100011101000111","0000111010101110101011101010","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111101011111010111110101","0000111111101111111011111110","0000111111001111110011111100","0000111110001111100011111000","0000111111111111111111111111","0000110000001100000011000000","0000000101010001010100010101","0001000000000000000000000000","0000001010100010101000101010","0000010001110100011101000111","0000110110101101101011011010","0000101011101010111010101110","0000111111111111111111111111","0000110011001100110011001100","0000101111111011111110111111","0000110010001100100011001000","0000111110111111101111111011","0000111000001110000011100000","0000110101011101010111010101","0000111111111111111111111111","0000101101001011010010110100","0000111010001110100011101000","0000111110111111101111111011","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111001101110011011100110","0000101101011011010110110101","0000111001101110011011100110","0000110000111100001111000011","0000010111100101111001011110","0000010100110101001101010011","0000000110000001100000011000","0001000000000000000000000000","0000011101000111010001110100","0000100001111000011110000111","0000100100011001000110010001","0000010111010101110101011101","0000000001100000011000000110","0000001110000011100000111000","0000001100010011000100110001","0000010001110100011101000111","0000011010100110101001101010","0000000001010000010100000101","0000101010111010101110101011","0000111010011110100111101001","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111100111111001111110011","0000111100011111000111110001","0000010000110100001101000011","0000000101110001011100010111","0000001001100010011000100110","0000011100010111000101110001","0000001000010010000100100001","0000001110110011101100111011","0000001100110011001100110011","0000101101001011010010110100","0000110101011101010111010101","0000010101010101010101010101","0000100100001001000010010000","0000101010011010100110101001","0000111111111111111111111111","0000111110111111101111111011","0000111101011111010111110101","0000111110101111101011111010","0000110111111101111111011111","0000101010001010100010101000","0000110101101101011011010110","0000101011011010110110101101","0000111010101110101011101010","0000110111011101110111011101","0000110001001100010011000100","0000100011101000111010001110","0000100101011001010110010101","0000100000111000001110000011","0000010010000100100001001000","0000011001110110011101100111","0000101110011011100110111001","0000110101111101011111010111","0000110110011101100111011001","0000110010001100100011001000","0000110000111100001111000011","0000011100100111001001110010","0000000010100000101000001010","0000000011010000110100001101","0000011011010110110101101101","0000100011001000110010001100","0000100111001001110010011100","0000011111110111111101111111","0000100001001000010010000100","0000010100100101001001010010","0000101100001011000010110000","0000011101110111011101110111","0000000010110000101100001011","0000110010111100101111001011","0000110000011100000111000001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111101101111011011110110","0000111010101110101011101010","0000111111111111111111111111","0000111110001111100011111000","0000111111111111111111111111","0000110000011100000111000001","0000001101100011011000110110","0000000001110000011100000111","0000000100100001001000010010","0000001110110011101100111011","0000100110111001101110011011","0000101001011010010110100101","0000101110011011100110111001","0000101101111011011110110111","0000101110001011100010111000","0000111000011110000111100001","0000111010011110100111101001","0000111010011110100111101001","0000111100111111001111110011","0000111011011110110111101101","0000101111011011110110111101","0000111111111111111111111111","0000111101001111010011110100","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000110110001101100011011000","0000111111111111111111111111","0000111001111110011111100111","0000011111000111110001111100","0000011111000111110001111100","0000011101110111011101110111","0000000010100000101000001010","0000000011100000111000001110","0000011111100111111001111110","0000101001011010010110100101","0000101111011011110110111101","0000110001101100011011000110","0000100011011000110110001101","0000000001100000011000000110","0000001110000011100000111000","0000011000010110000101100001","0000001110110011101100111011","0001000000000000000000000000","0000110111001101110011011100","0000111011111110111111101111","0000111111001111110011111100","0000111011101110111011101110","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000110101001101010011010100","0001000000000000000000000000","0001000000000000000000000000","0000010011100100111001001110","0000000111000001110000011100","0000001110100011101000111010","0000010101010101010101010101","0000011110000111100001111000","0000110110011101100111011001","0000011110110111101101111011","0000100100001001000010010000","0000100000101000001010000010","0000111100111111001111110011","0000110101111101011111010111","0000100110001001100010011000","0000100100011001000110010001","0000101010011010100110101001","0000101111111011111110111111","0000110111111101111111011111","0000101010101010101010101010","0000101011111010111110101111","0000101101001011010010110100","0000011111110111111101111111","0000011001000110010001100100","0000001100000011000000110000","0000010000000100000001000000","0000001100010011000100110001","0000010110000101100001011000","0000100100111001001110010011","0000101011011010110110101101","0000110001001100010011000100","0000110000101100001011000010","0000100100011001000110010001","0000001011100010111000101110","0000010010010100100101001001","0000000000100000001000000010","0000001011000010110000101100","0000001101000011010000110100","0000010110000101100001011000","0000011100110111001101110011","0000100110111001101110011011","0000100110111001101110011011","0000000111010001110100011101","0000000001110000011100000111","0000101100001011000010110000","0000110110101101101011011010","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111101111111011111110111","0000100110011001100110011001","0000000001000000010000000100","0000000010100000101000001010","0000011111100111111001111110","0000100111111001111110011111","0000011100000111000001110000","0000100010101000101010001010","0000101010001010100010101000","0000101001001010010010100100","0000101101001011010010110100","0000110011001100110011001100","0000110111111101111111011111","0000111110001111100011111000","0000111000101110001011100010","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111110111111101111111011","0000111101001111010011110100","0000100011011000110110001101","0000101001011010010110100101","0000100000101000001010000010","0000001111110011111100111111","0000000111110001111100011111","0000101011001010110010101100","0000111011011110110111101101","0000111111111111111111111111","0000111100011111000111110001","0000111101011111010111110101","0000100110111001101110011011","0000011001100110011001100110","0000001001010010010100100101","0000010001000100010001000100","0000010001000100010001000100","0000001001000010010000100100","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111110011111100111111001","0000111101111111011111110111","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000100010011000100110001001","0001000000000000000000000000","0001000000000000000000000000","0000001111000011110000111100","0000001100010011000100110001","0000001110000011100000111000","0000010110010101100101011001","0000100001001000010010000100","0000011011100110111001101110","0000100100101001001010010010","0000011100000111000001110000","0000101101111011011110110111","0000111010001110100011101000","0000111010001110100011101000","0000111001011110010111100101","0000110100101101001011010010","0000110100011101000111010001","0000110100101101001011010010","0000100111111001111110011111","0000101011001010110010101100","0000100011101000111010001110","0000010010100100101001001010","0000001010100010101000101010","0000011110010111100101111001","0000010011110100111101001111","0000011001110110011101100111","0000011000000110000001100000","0000010110000101100001011000","0000101000101010001010100010","0000110011111100111111001111","0000110001101100011011000110","0000100000011000000110000001","0000001111100011111000111110","0000010010010100100101001001","0000011011000110110001101100","0000001111010011110100111101","0000000011000000110000001100","0000001011010010110100101101","0000010111100101111001011110","0000001010010010100100101001","0000001101000011010000110100","0001000000000000000000000000","0000100001001000010010000100","0000111111011111110111111101","0000111010101110101011101010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111011011110110111101101","0000111010001110100011101000","0000111111111111111111111111","0000111111111111111111111111","0000110001101100011011000110","0000010000110100001101000011","0000000010100000101000001010","0000010000100100001001000010","0000011111000111110001111100","0000011100000111000001110000","0000011100000111000001110000","0000011010100110101001101010","0000010111000101110001011100","0000011010000110100001101000","0000101000011010000110100001","0000100111011001110110011101","0000110101101101011011010110","0000100100011001000110010001","0000111010011110100111101001","0000111100101111001011110010","0000111110101111101011111010","0000111110111111101111111011","0000111111001111110011111100","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000101111111011111110111111","0000111000011110000111100001","0000101001011010010110100101","0000010011110100111101001111","0000000001010000010100000101","0000110000001100000011000000","0000110000001100000011000000","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000100101011001010110010101","0000011110010111100101111001","0000001001000010010000100100","0000001011010010110100101101","0001000000000000000000000000","0000100101111001011110010111","0000111001001110010011100100","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111011001110110011101100","0000111111111111111111111111","0000111100011111000111110001","0000001101010011010100110101","0000000101000001010000010100","0000000101000001010000010100","0000010111000101110001011100","0000001110100011101000111010","0000001010000010100000101000","0000010101100101011001010110","0000001011000010110000101100","0000010110000101100001011000","0000100011111000111110001111","0000110001001100010011000100","0000111111111111111111111111","0000111111111111111111111111","0000111011001110110011101100","0000111010001110100011101000","0000110100111101001111010011","0000111000011110000111100001","0000101111111011111110111111","0000110000111100001111000011","0000100100001001000010010000","0000100010101000101010001010","0000100010101000101010001010","0000010010110100101101001011","0000101010011010100110101001","0000110011001100110011001100","0000010111100101111001011110","0000001110100011101000111010","0000101000011010000110100001","0000110101101101011011010110","0000110100001101000011010000","0000101000101010001010100010","0000011011000110110001101100","0000100010011000100110001001","0000100001001000010010000100","0000011011110110111101101111","0000010111000101110001011100","0000010100010101000101010001","0000011001010110010101100101","0000000001000000010000000100","0000001111110011111100111111","0000110010111100101111001011","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111110101111101011111010","0000111100011111000111110001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111101111111011111110111","0000111110111111101111111011","0000111110101111101011111010","0000111111001111110011111100","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000110101111101011111010111","0000011110010111100101111001","0001000000000000000000000000","0000000010100000101000001010","0000011000000110000001100000","0000001101110011011100110111","0000010011100100111001001110","0000001110100011101000111010","0000000101110001011100010111","0000001100000011000000110000","0000001111000011110000111100","0000010111110101111101011111","0000010110100101101001011010","0000100011111000111110001111","0000110011011100110111001101","0000111101001111010011110100","0000111011101110111011101110","0000111100001111000011110000","0000111111111111111111111111","0000111010101110101011101010","0000101111101011111010111110","0000101010111010101110101011","0000100001001000010010000100","0000001101000011010000110100","0001000000000000000000000000","0000101110001011100010111000","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000110010111100101111001011","0000101111011011110110111101","0000010110100101101001011010","0000010101010101010101010101","0000001000110010001100100011","0000000011110000111100001111","0000101011111010111110101111","0000110111011101110111011101","0000111110111111101111111011","0000111111111111111111111111","0000111110011111100111111001","0000111110101111101011111010","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000010000010100000101000001","0000000000100000001000000010","0000001000010010000100100001","0000010010110100101101001011","0000000000110000001100000011","0000001111100011111000111110","0000010100010101000101010001","0000001111110011111100111111","0000010000100100001001000010","0000011000010110000101100001","0000101011111010111110101111","0000101011001010110010101100","0000101110111011101110111011","0000011100110111001101110011","0000010110000101100001011000","0000001101010011010100110101","0000001100100011001000110010","0000000101110001011100010111","0000001101110011011100110111","0000010001000100010001000100","0000010000010100000101000001","0000010110010101100101011001","0000001110110011101100111011","0000001100110011001100110011","0000001101100011011000110110","0000001001100010011000100110","0000011101000111010001110100","0000110101111101011111010111","0000101100011011000110110001","0000100001011000010110000101","0000110101101101011011010110","0000111011001110110011101100","0000110011101100111011001110","0000101000001010000010100000","0000100011001000110010001100","0000010111000101110001011100","0000000101000001010000010100","0000100110101001101010011010","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111100111111001111110011","0000111111111111111111111111","0000111110001111100011111000","0000111100101111001011110010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111101011111010111110101","0000111101111111011111110111","0000111111111111111111111111","0000111111101111111011111110","0000110010001100100011001000","0000011011010110110101101101","0000001000110010001100100011","0000000111010001110100011101","0000010111100101111001011110","0000010011010100110101001101","0000001010110010101100101011","0000001110000011100000111000","0000001000000010000000100000","0000000010000000100000001000","0000001001110010011100100111","0000011000100110001001100010","0000010100100101001001010010","0000010101010101010101010101","0000100001001000010010000100","0000100110001001100010011000","0000101011101010111010101110","0000100011111000111110001111","0000011010000110100001101000","0000001111010011110100111101","0000000000100000001000000010","0000010101110101011101010111","0000110101101101011011010110","0000111111101111111011111110","0000111110101111101011111010","0000111100101111001011110010","0000111111111111111111111111","0000111111101111111011111110","0000111011011110110111101101","0000100110101001101010011010","0000101001111010011110100111","0000011000100110001001100010","0000001110110011101100111011","0000000101010001010100010101","0000011001110110011101100111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111011111110111111101","0000111010011110100111101001","0000100010001000100010001000","0000000101100001011000010110","0001000000000000000000000000","0000001010000010100000101000","0000001100110011001100110011","0000000110010001100100011001","0000000001110000011100000111","0000000111010001110100011101","0001000000000000000000000000","0000000100000001000000010000","0000001100110011001100110011","0000001101000011010000110100","0000010011110100111101001111","0000011111100111111001111110","0000101011101010111010101110","0000110011101100111011001110","0000110101101101011011010110","0000111010001110100011101000","0000111101011111010111110101","0000111111111111111111111111","0000111010111110101111101011","0000110000001100000011000000","0000100010011000100110001001","0000011000100110001001100010","0000010100110101001101010011","0000011100010111000101110001","0000100101101001011010010110","0000100100001001000010010000","0000101101111011011110110111","0000111010111110101111101011","0000111111111111111111111111","0000111110001111100011111000","0000101111001011110010111100","0000001111100011111000111110","0000001110110011101100111011","0000110001011100010111000101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111101101111011011110110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111001001110010011100100","0000110010111100101111001011","0000100101111001011110010111","0001000000000000000000000000","0000011100000111000001110000","0000100001111000011110000111","0000010110100101101001011010","0000100011001000110010001100","0000010111110101111101011111","0000011001010110010101100101","0000000111000001110000011100","0000001010010010100100101001","0000011001100110011001100110","0000011111110111111101111111","0000011110010111100101111001","0000010100110101001101010011","0000001100010011000100110001","0001000000000000000000000000","0000001110010011100100111001","0000110000101100001011000010","0000111111011111110111111101","0000111110011111100111111001","0000111111111111111111111111","0000111110001111100011111000","0000110111011101110111011101","0000111010001110100011101000","0000110010011100100111001001","0000101011001010110010101100","0000010100100101001001010010","0000010110000101100001011000","0000011100100111001001110010","0000010101100101011001010110","0000000010100000101000001010","0000110011001100110011001100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000101011101010111010101110","0000010010110100101101001011","0000000001000000010000000100","0000001100110011001100110011","0000100101001001010010010100","0000011100110111001101110011","0000010110000101100001011000","0000001001110010011100100111","0001000000000000000000000000","0000101000001010000010100000","0000111011111110111111101111","0000111110011111100111111001","0000111110101111101011111010","0000111111111111111111111111","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111010101110101011101010","0000101000111010001110100011","0000101010101010101010101010","0000011110010111100101111001","0000010111010101110101011101","0000100111001001110010011100","0000101000011010000110100001","0000100001011000010110000101","0000110010111100101111001011","0000111111111111111111111111","0000111001001110010011100100","0000101000011010000110100001","0000001011000010110000101100","0000000001000000010000000100","0000100101011001010110010101","0000111111111111111111111111","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111001111110011111100","0000111110111111101111111011","0000111110111111101111111011","0000111111001111110011111100","0000111111001111110011111100","0000111110111111101111111011","0000111110101111101011111010","0000111001111110011111100111","0000010010010100100101001001","0000001101010011010100110101","0000011101000111010001110100","0000011110100111101001111010","0000100010001000100010001000","0000010101010101010101010101","0000010110010101100101011001","0000010100010101000101010001","0000001100000011000000110000","0000000011110000111100001111","0000001100100011001000110010","0000010001110100011101000111","0000100011001000110010001100","0000110111101101111011011110","0000111100101111001011110010","0000111111111111111111111111","0000111100101111001011110010","0000111101011111010111110101","0000111111111111111111111111","0000111111001111110011111100","0000111100001111000011110000","0000110100101101001011010010","0000100111001001110010011100","0000001111110011111100111111","0000100110001001100010011000","0000101011011010110110101101","0000101011011010110110101101","0000000111100001111000011110","0000010110010101100101011001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000110011001100110011001100","0000100001111000011110000111","0000000001110000011100000111","0000000101100001011000010110","0000011010110110101101101011","0000010111100101111001011110","0000010100100101001001010010","0000010110110101101101011011","0000010111100101111001011110","0000011010010110100101101001","0000101101101011011010110110","0000111000011110000111100001","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110000001100000011000000","0000100011101000111010001110","0000101011101010111010101110","0000100001001000010010000100","0000101010001010100010101000","0000111001001110010011100100","0000101101111011011110110111","0000101100001011000010110000","0000110100101101001011010010","0000100001001000010010000100","0000011100010111000101110001","0000000000010000000100000001","0000000110110001101100011011","0000101011111010111110101111","0000111110111111101111111011","0000111110101111101011111010","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111011111110111111101","0000111111101111111011111110","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000110100001101000011010000","0000011001000110010001100100","0000000100110001001100010011","0000010000100100001001000010","0000101011001010110010101100","0000101100101011001010110010","0000011110000111100001111000","0000010011000100110001001100","0000011000100110001001100010","0000011001110110011101100111","0000100001101000011010000110","0000101011001010110010101100","0000110110101101101011011010","0000111110111111101111111011","0000111100001111000011110000","0000111110101111101011111010","0000111111011111110111111101","0000110111011101110111011101","0000111010101110101011101010","0000111110011111100111111001","0000101110011011100110111001","0000100000101000001010000010","0000110011011100110111001101","0000101101101011011010110110","0000111101101111011011110110","0000100001111000011110000111","0000000100100001001000010010","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111111111111111111111","0000111110101111101011111010","0000111100001111000011110000","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000110100101101001011010010","0000010011010100110101001101","0001000000000000000000000000","0000100110011001100110011001","0000101100001011000010110000","0000011011110110111101101111","0000100011011000110110001101","0000100010111000101110001011","0000011111010111110101111101","0000011010010110100101101001","0000100100011001000110010001","0000101101101011011010110110","0000111000111110001111100011","0000110000111100001111000011","0000110100101101001011010010","0000111000001110000011100000","0000011111000111110001111100","0000100111111001111110011111","0000110101111101011111010111","0000101101111011011110110111","0000100000011000000110000001","0000010100010101000101010001","0000000010100000101000001010","0001000000000000000000000000","0000010110000101100001011000","0000110011011100110111001101","0000111111111111111111111111","0000111100101111001011110010","0000111111011111110111111101","0000111111111111111111111111","0000111111001111110011111100","0000111110111111101111111011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111011111110111111101","0000111111001111110011111100","0000111110111111101111111011","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111110011111100111111001","0000111101111111011111110111","0000111111111111111111111111","0000110101011101010111010101","0000011011010110110101101101","0000000001100000011000000110","0000010000000100000001000000","0000100001111000011110000111","0000100100001001000010010000","0000101001011010010110100101","0000110010111100101111001011","0000110001101100011011000110","0000011111110111111101111111","0000011011100110111001101110","0000101110011011100110111001","0000110011011100110111001101","0000110110111101101111011011","0000110010111100101111001011","0000110101011101010111010101","0000111000111110001111100011","0000101101101011011010110110","0000100010111000101110001011","0000110001101100011011000110","0000110010001100100011001000","0000111100001111000011110000","0000101000111010001110100011","0000000010100000101000001010","0000101101011011010110110101","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111101111111011111110111","0000111101101111011011110110","0000111100111111001111110011","0000111111101111111011111110","0000101011001010110010101100","0000001110000011100000111000","0001000000000000000000000000","0000001100000011000000110000","0000010011010100110101001101","0000011000010110000101100001","0000010111010101110101011101","0000011110000111100001111000","0000011001110110011101100111","0000011010010110100101101001","0000011001100110011001100110","0000101000001010000010100000","0000100100111001001110010011","0000011111100111111001111110","0000010101000101010001010100","0000010100100101001001010010","0000000001110000011100000111","0001000000000000000000000000","0000001110010011100100111001","0000011101000111010001110100","0000110000111100001111000011","0000111001001110010011100100","0000111001011110010111100101","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111100101111001011110010","0000111100111111001111110011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110011111100111111001","0000111101111111011111110111","0000111101111111011111110111","0000111110001111100011111000","0000111101101111011011110110","0000111101011111010111110101","0000111110111111101111111011","0000111111111111111111111111","0000111110111111101111111011","0000111110101111101011111010","0000111100011111000111110001","0000111110011111100111111001","0000111111111111111111111111","0000110101111101011111010111","0000100000011000000110000001","0000001110100011101000111010","0000001100110011001100110011","0000010110100101101001011010","0000100011001000110010001100","0000100110101001101010011010","0000110001001100010011000100","0000110110101101101011011010","0000101011001010110010101100","0000101101101011011010110110","0000101110111011101110111011","0000100111011001110110011101","0000100101011001010110010101","0000100001101000011010000110","0000011101110111011101110111","0000101011001010110010101100","0000101100011011000110110001","0000110100111101001111010011","0000101010111010101110101011","0001000000000000000000000000","0000110000101100001011000010","0000111111111111111111111111","0000111010101110101011101010","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111110111111101111111011","0000111111111111111111111111","0000111111001111110011111100","0000111100111111001111110011","0000111111111111111111111111","0000111101111111011111110111","0000111111111111111111111111","0000111101011111010111110101","0000110101001101010011010100","0000100001101000011010000110","0000010100100101001001010010","0000001100000011000000110000","0000000111110001111100011111","0001000000000000000000000000","0000000000100000001000000010","0001000000000000000000000000","0000000010100000101000001010","0001000000000000000000000000","0000000101000001010000010100","0000001011100010111000101110","0000010110100101101001011010","0000011110010111100101111001","0000101101101011011010110110","0000110100011101000111010001","0000111011111110111111101111","0000111110011111100111111001","0000111010101110101011101010","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111010111110101111101011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111101111111011111110","0000111111101111111011111110","0000111110111111101111111011","0000111111111111111111111111","0000111011011110110111101101","0000111110111111101111111011","0000111111011111110111111101","0000111110111111101111111011","0000111111111111111111111111","0000111100101111001011110010","0000111100101111001011110010","0000111111111111111111111111","0000110100011101000111010001","0000010110110101101101011011","0000001101010011010100110101","0000010010100100101001001010","0000011110010111100101111001","0000100000011000000110000001","0000101000011010000110100001","0000101001001010010010100100","0000101011101010111010101110","0000100111111001111110011111","0000100001001000010010000100","0000100001001000010010000100","0000100101101001011010010110","0000101010001010100010101000","0000110001011100010111000101","0000010111100101111001011110","0000000011100000111000001110","0000110010111100101111001011","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111011111110111111101111","0000111111101111111011111110","0000111111111111111111111111","0000111111011111110111111101","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111101001111010011110100","0000111101001111010011110100","0000111111111111111111111111","0000110110111101101111011011","0000110110011101100111011001","0000110111101101111011011110","0000110110111101101111011011","0000111001011110010111100101","0000110010101100101011001010","0000110001101100011011000110","0000110001101100011011000110","0000110111111101111111011111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111110111111101111111011","0000111011011110110111101101","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111011001110110011101100","0000111101001111010011110100","0000111111111111111111111111","0000111110011111100111111001","0000111100111111001111110011","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111100011111000111110001","0000111011001110110011101100","0000111100111111001111110011","0000111110111111101111111011","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111101011111010111110101","0000111111111111111111111111","0000111111111111111111111111","0000111101111111011111110111","0000111101011111010111110101","0000111111111111111111111111","0000111010111110101111101011","0000110110001101100011011000","0000100010101000101010001010","0000001100110011001100110011","0000000110100001101000011010","0000001000100010001000100010","0000001100000011000000110000","0000010111000101110001011100","0000010110010101100101011001","0000001110000011100000111000","0000010001010100010101000101","0000010011000100110001001100","0000000010100000101000001010","0000011000110110001101100011","0000111001101110011011100110","0000111010101110101011101010","0000111111111111111111111111","0000111111101111111011111110","0000111110011111100111111001","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111101101111011011110110","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111110011111100111111001","0000111111011111110111111101","0000111111111111111111111111","0000111111111111111111111111","0000111111001111110011111100","0000111111101111111011111110","0000111110001111100011111000","0000111111111111111111111111","0000111101011111010111110101","0000111111011111110111111101","0000111111111111111111111111","0000111110001111100011111000","0000111110011111100111111001","0000111111101111111011111110","0000111111111111111111111111","0000111111101111111011111110","0000111110111111101111111011","0000111110001111100011111000","0000111110101111101011111010","0000111110001111100011111000","0000111111111111111111111111","0000111111011111110111111101","0000111110001111100011111000","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111110001111100011111000","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111100001111000011110000","0000111101101111011011110110","0000111111111111111111111111","0000111101101111011011110110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111",
		"0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111000011110000111100001","0000110001011100010111000101","0000100111011001110110011101","0000011101110111011101110111","0000010111000101110001011100","0000011000000110000001100000","0000100001101000011010000110","0000101011101010111010101110","0000111001011110010111100101","0000111111001111110011111100","0000111111111111111111111111","0000111110101111101011111010","0000111111111111111111111111","0000111111111111111111111111","0000111110111111101111111011","0000111111101111111011111110","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111","0000111111111111111111111111"

	);
begin
	process (clk)
	begin
		if rising_edge(clk) then
			if en = '1' then
				if addr <= "1100010001111010" then --1100010001111001
					data <= ROM(TO_INTEGER(addr)); 
				else
					data <= "0001000000000000000000000000"; 
				end if;
			else
				data <= "0001000000000000000000000000"; 
			end if;
		end if;
	end process;
end imp;